LIBRARY ieee;
USE ieee.std_logic_1164.all; 
use ieee.std_logic_unsigned.all;

LIBRARY work;

ENTITY VGA_REGS IS 
	PORT
	(
		CLK     : IN  STD_LOGIC;
		RESET_n : IN  STD_LOGIC;

--		CSmem   : IN  STD_LOGIC;
		CSreg   : IN  STD_LOGIC;
		A       : IN  STD_LOGIC_VECTOR(16 DOWNTO 0);
		D       : IN  STD_LOGIC_VECTOR(7 DOWNTO 0);

		CONTROL : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
--		CONTROLx: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		HSCROLL : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		VSCROLL : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);

		HCURSOR : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		VCURSOR : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);

		VDo     : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		VA      : OUT STD_LOGIC_VECTOR(16 DOWNTO 0);
		VWE     : OUT STD_LOGIC;
		BLE     : OUT STD_LOGIC;
		BHE     : OUT STD_LOGIC
	);
END VGA_REGS;

ARCHITECTURE bdf_type OF VGA_REGS IS 

SIGNAL	REG0       :  STD_LOGIC;
SIGNAL	REG00      :  STD_LOGIC;
SIGNAL	REG01      :  STD_LOGIC;
SIGNAL	REG02      :  STD_LOGIC;
SIGNAL	REG1       :  STD_LOGIC;
SIGNAL	REG2       :  STD_LOGIC;
SIGNAL	REG3       :  STD_LOGIC;
SIGNAL	REG4       :  STD_LOGIC;
SIGNAL	REG40      :  STD_LOGIC;
SIGNAL	REG41      :  STD_LOGIC;
SIGNAL	REG5       :  STD_LOGIC;
SIGNAL	REG6       :  STD_LOGIC;
SIGNAL	REG7       :  STD_LOGIC;

SIGNAL	REG_ADDR    : STD_LOGIC_VECTOR(17 DOWNTO 0);
SIGNAL	REG_DATA    : STD_LOGIC_VECTOR(7 DOWNTO 0);
--SIGNAL	REG_ACCCTRL : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	REG_CTRL    : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	REG_HSCROLL : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	REG_VSCROLL : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	REG_COLOR   : STD_LOGIC_VECTOR(15 DOWNTO 0);
--SIGNAL	REG_CTRLx   : STD_LOGIC_VECTOR(7 DOWNTO 0);
--SIGNAL	REG_ABUF    : STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	REG_INC     : STD_LOGIC_VECTOR(5 DOWNTO 0);

SIGNAL	BHiEn :  STD_LOGIC;
SIGNAL	BLoEn :  STD_LOGIC;

SIGNAL	WRCPU  :  STD_LOGIC;

BEGIN
-------------------------------------------------------------------------------
-- REGISTERS
-------------------------------------------------------------------------------
REG0 <= NOT(CSreg) AND NOT(A(2)) AND NOT(A(1)) AND NOT(A(0));
REG1 <= NOT(CSreg) AND NOT(A(2)) AND NOT(A(1)) AND     A(0);
REG2 <= NOT(CSreg) AND NOT(A(2)) AND     A(1)  AND NOT(A(0));
REG3 <= NOT(CSreg) AND NOT(A(2)) AND     A(1)  AND     A(0);
REG4 <= NOT(CSreg) AND     A(2)  AND NOT(A(1)) AND NOT(A(0));
REG5 <= NOT(CSreg) AND     A(2)  AND NOT(A(1)) AND     A(0);
REG6 <= NOT(CSreg) AND     A(2)  AND     A(1)  AND NOT(A(0));
REG7 <= NOT(CSreg) AND     A(2)  AND     A(1)  AND     A(0);

--REG00 <= REG0 AND NOT(REG_ABUF(1)) AND NOT(REG_ABUF(0));
--REG01 <= REG0 AND NOT(REG_ABUF(1)) AND     REG_ABUF(0) ;
--REG02 <= REG0 AND     REG_ABUF(1)  AND NOT(REG_ABUF(0));

--REG40 <= REG4 AND NOT(REG_ABUF(0));
--REG41 <= REG4 AND     REG_ABUF(0) ;

PROCESS(RESET_n, REG7, CLK)
BEGIN
  IF (RESET_n = '0') THEN
    CONTROL  <= (OTHERS => '0');
--    CONTROLx <= "00000000";
  ELSIF (RISING_EDGE(REG7)) THEN
--    IF (D(7) = '0' ) THEN
      CONTROL  <= D(7 DOWNTO 0);
--    ELSE
--      CONTROLx <= D(6 DOWNTO 0);
--    END IF;
  END IF;
END PROCESS;

PROCESS(RESET_n, REG6, CLK)
BEGIN
  IF (RESET_n = '0') THEN
    VSCROLL <= (OTHERS => '0');
  ELSIF (RISING_EDGE(REG6)) THEN
    VSCROLL <= D;
  END IF;
END PROCESS;

PROCESS(RESET_n, REG5, CLK)
BEGIN
  IF (RESET_n = '0') THEN
    HSCROLL <= (OTHERS => '0');
  ELSIF (RISING_EDGE(REG5)) THEN
    HSCROLL <= D;
  END IF;
END PROCESS;

PROCESS(RESET_n, REG4, CLK)
BEGIN
  IF (RESET_n = '0') THEN
    REG_COLOR( 7 DOWNTO  0) <= (OTHERS => '0');
  ELSIF (RISING_EDGE(REG4)) THEN
    REG_COLOR( 7 DOWNTO  0) <= D;
  END IF;
END PROCESS;

PROCESS(RESET_n, REG3, CLK)
BEGIN
  IF (RESET_n = '0') THEN
    VCURSOR <= (OTHERS => '0');
  ELSIF (RISING_EDGE(REG3)) THEN
    VCURSOR <= D(7 DOWNTO 0);
  END IF;
END PROCESS;

PROCESS(RESET_n, REG2, CLK)
BEGIN
  IF (RESET_n = '0') THEN
    HCURSOR <= (OTHERS => '0');
  ELSIF (RISING_EDGE(REG2)) THEN
    HCURSOR <= D(7 DOWNTO 0);
  END IF;
END PROCESS;

PROCESS(RESET_n, REG1, CLK)
BEGIN
  IF (RESET_n = '0') THEN
    REG_DATA <= (OTHERS => '0');
  ELSIF (RISING_EDGE(REG1)) THEN
    REG_DATA <= D;
--    REG_ADDR <= REG_ADDR + REG_INC;
  END IF;
END PROCESS;

PROCESS(RESET_n, REG0, CLK)
BEGIN
  IF (RESET_n = '0') THEN
    REG_ADDR( 5 DOWNTO  0) <= (OTHERS => '0');
    REG_ADDR(11 DOWNTO  6) <= (OTHERS => '0');
    REG_ADDR(17 DOWNTO 12) <= (OTHERS => '0');
    REG_INC <= (OTHERS => '0');
  ELSIF (RISING_EDGE(REG0)) THEN
    CASE D(7 DOWNTO 6) IS
    WHEN "00" => REG_ADDR( 5 DOWNTO  0) <= D( 5 DOWNTO  0);
    WHEN "01" => REG_ADDR(11 DOWNTO  6) <= D( 5 DOWNTO  0);
    WHEN "10" => REG_ADDR(17 DOWNTO 12) <= D( 5 DOWNTO  0);
    WHEN "11" => REG_INC <= D(5 DOWNTO  0);
    END CASE;
  END IF;
END PROCESS;

VA    <= REG_ADDR(17 DOWNTO 1);
VDo   <= REG_DATA;
BLE   <= REG_ADDR(0);
BHE   <= NOT(REG_ADDR(0));
VWE   <= NOT(REG1);
-------------------------------------------------------------------------------
END bdf_type;
