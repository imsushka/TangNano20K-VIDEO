LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY count IS 
	PORT
	(
		CLK :   IN  STD_LOGIC;
		SClr :  IN  STD_LOGIC; -- 0 reset / 1 count
		Q :     OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
	);
END count;

ARCHITECTURE bdf_type OF count IS 

SIGNAL	D :  STD_LOGIC_VECTOR(11 DOWNTO 0);
SIGNAL	Q_SYNTH :  STD_LOGIC_VECTOR(11 DOWNTO 0);
SIGNAL	WIRE_0 :  STD_LOGIC;
SIGNAL	WIRE_1 :  STD_LOGIC;
SIGNAL	WIRE_2 :  STD_LOGIC;
SIGNAL	WIRE_3 :  STD_LOGIC;
SIGNAL	WIRE_4 :  STD_LOGIC;
SIGNAL	WIRE_5 :  STD_LOGIC;
SIGNAL	WIRE_6 :  STD_LOGIC;
SIGNAL	WIRE_7 :  STD_LOGIC;
SIGNAL	WIRE_8 :  STD_LOGIC;
SIGNAL	WIRE_9 :  STD_LOGIC;
SIGNAL	WIRE_10 :  STD_LOGIC;
SIGNAL	WIRE_11 :  STD_LOGIC;

SIGNAL	WIRE_00 :  STD_LOGIC;
SIGNAL	WIRE_01 :  STD_LOGIC;
SIGNAL	WIRE_02 :  STD_LOGIC;
SIGNAL	WIRE_03 :  STD_LOGIC;
SIGNAL	WIRE_04 :  STD_LOGIC;
SIGNAL	WIRE_05 :  STD_LOGIC;
SIGNAL	WIRE_06 :  STD_LOGIC;
SIGNAL	WIRE_07 :  STD_LOGIC;
SIGNAL	WIRE_08 :  STD_LOGIC;
SIGNAL	WIRE_09 :  STD_LOGIC;

BEGIN 

PROCESS(CLK)
BEGIN
IF (RISING_EDGE(CLK)) THEN
	Q_SYNTH(11 DOWNTO 0) <= D(11 DOWNTO 0);
END IF;
END PROCESS;

WIRE_0 <= NOT(Q_SYNTH(0));
D(0) <= SClr AND WIRE_0;

WIRE_1 <= Q_SYNTH(0) XOR Q_SYNTH(1);
D(1) <= SClr AND WIRE_1;

WIRE_01 <= Q_SYNTH(0) AND Q_SYNTH(1);
WIRE_2 <= Q_SYNTH(2) XOR WIRE_01;
D(2) <= SClr AND WIRE_2;

WIRE_02 <= WIRE_01 AND Q_SYNTH(2);
WIRE_3 <= Q_SYNTH(3) XOR WIRE_02;
D(3) <= SClr AND WIRE_3;

WIRE_03 <= WIRE_02 AND Q_SYNTH(3);
WIRE_4 <= Q_SYNTH(4) XOR WIRE_03;
D(4) <= SClr AND WIRE_4;

WIRE_04 <= WIRE_03 AND Q_SYNTH(4);
WIRE_5 <= Q_SYNTH(5) XOR WIRE_04;
D(5) <= SClr AND WIRE_5;

WIRE_05 <= WIRE_04 AND Q_SYNTH(5);
WIRE_6 <= Q_SYNTH(6) XOR WIRE_05;
D(6) <= SClr AND WIRE_6;

WIRE_06 <= WIRE_05 AND Q_SYNTH(6);
WIRE_7 <= Q_SYNTH(7) XOR WIRE_06;
D(7) <= SClr AND WIRE_7;

WIRE_07 <= WIRE_06 AND Q_SYNTH(7);
WIRE_8 <= Q_SYNTH(8) XOR WIRE_07;
D(8) <= SClr AND WIRE_8;

WIRE_08 <= WIRE_07 AND Q_SYNTH(8);
WIRE_9 <= Q_SYNTH(9) XOR WIRE_08;
D(9) <= SClr AND WIRE_9;

WIRE_09 <= WIRE_08 AND Q_SYNTH(9);
WIRE_10 <= Q_SYNTH(10) XOR WIRE_09;
D(10) <= SClr AND WIRE_10;

WIRE_00 <= WIRE_09 AND Q_SYNTH(10);
WIRE_11 <= Q_SYNTH(11) XOR WIRE_00;
D(11) <= SClr AND WIRE_11;

Q <= Q_SYNTH;

END bdf_type;