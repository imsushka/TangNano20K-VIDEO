library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
library work;

entity Video_Ram is
	port(
		clk    : in std_logic;

		addr_w : in std_logic_vector(15 downto 0);
		data_w : in std_logic_vector(15 downto 0);
		we     : in std_logic;
		le     : in std_logic;
		he     : in std_logic;

		addr_r : in std_logic_vector(15 downto 0);
		data_r : out std_logic_vector(15 downto 0)
	);
end Video_Ram;

architecture Behavioral of Video_Ram is
   
	constant ADDR_WIDTH : integer := 13;
	
	type ram_type is array (0 to 16383) of std_logic_vector(7 downto 0);
    
	-- ROM definition
	signal RAM_SCREEN_Lo: ram_type := (   -- 2^13-by-16
x"00",x"01",x"02",x"03",x"04",x"05",x"06",x"07",x"08",x"09",x"0A",x"0B",x"0C",x"0D",x"0E",x"0F",
x"10",x"11",x"12",x"13",x"14",x"15",x"16",x"17",x"18",x"19",x"1A",x"1B",x"1C",x"1D",x"1E",x"1F",
x"20",x"21",x"22",x"23",x"24",x"25",x"26",x"27",x"28",x"29",x"2A",x"2B",x"2C",x"2D",x"2E",x"2F",
x"30",x"31",x"32",x"33",x"34",x"35",x"36",x"37",x"38",x"39",x"3A",x"3B",x"3C",x"3D",x"3E",x"3F",
x"40",x"41",x"42",x"43",x"44",x"45",x"46",x"47",x"48",x"49",x"4A",x"4B",x"4C",x"4D",x"4E",x"4F",
x"50",x"51",x"52",x"53",x"54",x"55",x"56",x"57",x"58",x"59",x"5A",x"5B",x"5C",x"5D",x"5E",x"5F",
x"60",x"61",x"62",x"63",x"64",x"65",x"66",x"67",x"68",x"69",x"6A",x"6B",x"6C",x"6D",x"6E",x"6F",
x"70",x"71",x"72",x"73",x"74",x"75",x"76",x"77",x"78",x"79",x"7A",x"7B",x"7C",x"7D",x"7E",x"7F",
x"00",x"01",x"02",x"03",x"04",x"05",x"06",x"07",x"08",x"09",x"0A",x"0B",x"0C",x"0D",x"0E",x"0F",
x"10",x"11",x"12",x"13",x"14",x"15",x"16",x"17",x"18",x"19",x"1A",x"1B",x"1C",x"1D",x"1E",x"1F",
x"20",x"21",x"22",x"23",x"24",x"25",x"26",x"27",x"28",x"29",x"2A",x"2B",x"2C",x"2D",x"2E",x"2F",
x"30",x"31",x"32",x"33",x"34",x"35",x"36",x"37",x"38",x"39",x"3A",x"3B",x"3C",x"3D",x"3E",x"3F",
x"40",x"41",x"42",x"43",x"44",x"45",x"46",x"47",x"48",x"49",x"4A",x"4B",x"4C",x"4D",x"4E",x"4F",
x"50",x"51",x"52",x"53",x"54",x"55",x"56",x"57",x"58",x"59",x"5A",x"5B",x"5C",x"5D",x"5E",x"5F",
x"60",x"61",x"62",x"63",x"64",x"65",x"66",x"67",x"68",x"69",x"6A",x"6B",x"6C",x"6D",x"6E",x"6F",
x"70",x"71",x"72",x"73",x"74",x"75",x"76",x"77",x"78",x"79",x"7A",x"7B",x"7C",x"7D",x"7E",x"7F",

x"00",x"01",x"02",x"03",x"04",x"05",x"06",x"07",x"08",x"09",x"0A",x"0B",x"0C",x"0D",x"0E",x"0F",
x"10",x"11",x"12",x"13",x"14",x"15",x"16",x"17",x"18",x"19",x"1A",x"1B",x"1C",x"1D",x"1E",x"1F",
x"20",x"21",x"22",x"23",x"24",x"25",x"26",x"27",x"28",x"29",x"2A",x"2B",x"2C",x"2D",x"2E",x"2F",
x"30",x"31",x"32",x"33",x"34",x"35",x"36",x"37",x"38",x"39",x"3A",x"3B",x"3C",x"3D",x"3E",x"3F",
x"40",x"41",x"42",x"43",x"44",x"45",x"46",x"47",x"48",x"49",x"4A",x"4B",x"4C",x"4D",x"4E",x"4F",
x"50",x"51",x"52",x"53",x"54",x"55",x"56",x"57",x"58",x"59",x"5A",x"5B",x"5C",x"5D",x"5E",x"5F",
x"60",x"61",x"62",x"63",x"64",x"65",x"66",x"67",x"68",x"69",x"6A",x"6B",x"6C",x"6D",x"6E",x"6F",
x"70",x"71",x"72",x"73",x"74",x"75",x"76",x"77",x"78",x"79",x"7A",x"7B",x"7C",x"7D",x"7E",x"7F",
x"00",x"01",x"02",x"03",x"04",x"05",x"06",x"07",x"08",x"09",x"0A",x"0B",x"0C",x"0D",x"0E",x"0F",
x"10",x"11",x"12",x"13",x"14",x"15",x"16",x"17",x"18",x"19",x"1A",x"1B",x"1C",x"1D",x"1E",x"1F",
x"20",x"21",x"22",x"23",x"24",x"25",x"26",x"27",x"28",x"29",x"2A",x"2B",x"2C",x"2D",x"2E",x"2F",
x"30",x"31",x"32",x"33",x"34",x"35",x"36",x"37",x"38",x"39",x"3A",x"3B",x"3C",x"3D",x"3E",x"3F",
x"40",x"41",x"42",x"43",x"44",x"45",x"46",x"47",x"48",x"49",x"4A",x"4B",x"4C",x"4D",x"4E",x"4F",
x"50",x"51",x"52",x"53",x"54",x"55",x"56",x"57",x"58",x"59",x"5A",x"5B",x"5C",x"5D",x"5E",x"5F",
x"60",x"61",x"62",x"63",x"64",x"65",x"66",x"67",x"68",x"69",x"6A",x"6B",x"6C",x"6D",x"6E",x"6F",
x"70",x"71",x"72",x"73",x"74",x"75",x"76",x"77",x"78",x"79",x"7A",x"7B",x"7C",x"7D",x"7E",x"7F",

x"00",x"01",x"02",x"03",x"04",x"05",x"06",x"07",x"08",x"09",x"0A",x"0B",x"0C",x"0D",x"0E",x"0F",
x"10",x"11",x"12",x"13",x"14",x"15",x"16",x"17",x"18",x"19",x"1A",x"1B",x"1C",x"1D",x"1E",x"1F",
x"20",x"21",x"22",x"23",x"24",x"25",x"26",x"27",x"28",x"29",x"2A",x"2B",x"2C",x"2D",x"2E",x"2F",
x"30",x"31",x"32",x"33",x"34",x"35",x"36",x"37",x"38",x"39",x"3A",x"3B",x"3C",x"3D",x"3E",x"3F",
x"40",x"41",x"42",x"43",x"44",x"45",x"46",x"47",x"48",x"49",x"4A",x"4B",x"4C",x"4D",x"4E",x"4F",
x"50",x"51",x"52",x"53",x"54",x"55",x"56",x"57",x"58",x"59",x"5A",x"5B",x"5C",x"5D",x"5E",x"5F",
x"60",x"61",x"62",x"63",x"64",x"65",x"66",x"67",x"68",x"69",x"6A",x"6B",x"6C",x"6D",x"6E",x"6F",
x"70",x"71",x"72",x"73",x"74",x"75",x"76",x"77",x"78",x"79",x"7A",x"7B",x"7C",x"7D",x"7E",x"7F",
x"00",x"01",x"02",x"03",x"04",x"05",x"06",x"07",x"08",x"09",x"0A",x"0B",x"0C",x"0D",x"0E",x"0F",
x"10",x"11",x"12",x"13",x"14",x"15",x"16",x"17",x"18",x"19",x"1A",x"1B",x"1C",x"1D",x"1E",x"1F",
x"20",x"21",x"22",x"23",x"24",x"25",x"26",x"27",x"28",x"29",x"2A",x"2B",x"2C",x"2D",x"2E",x"2F",
x"30",x"31",x"32",x"33",x"34",x"35",x"36",x"37",x"38",x"39",x"3A",x"3B",x"3C",x"3D",x"3E",x"3F",
x"40",x"41",x"42",x"43",x"44",x"45",x"46",x"47",x"48",x"49",x"4A",x"4B",x"4C",x"4D",x"4E",x"4F",
x"50",x"51",x"52",x"53",x"54",x"55",x"56",x"57",x"58",x"59",x"5A",x"5B",x"5C",x"5D",x"5E",x"5F",
x"60",x"61",x"62",x"63",x"64",x"65",x"66",x"67",x"68",x"69",x"6A",x"6B",x"6C",x"6D",x"6E",x"6F",
x"70",x"71",x"72",x"73",x"74",x"75",x"76",x"77",x"78",x"79",x"7A",x"7B",x"7C",x"7D",x"7E",x"7F",

x"00",x"01",x"02",x"03",x"04",x"05",x"06",x"07",x"08",x"09",x"0A",x"0B",x"0C",x"0D",x"0E",x"0F",
x"20",x"20",x"20",x"20",x"53",x"55",x"48",x"41",x"53",x"48",x"4B",x"41",x"20",x"20",x"20",x"20",
x"53",x"56",x"49",x"4E",x"20",x"20",x"20",x"20",x"28",x"29",x"2A",x"2B",x"2C",x"2D",x"2E",x"2F",
x"30",x"31",x"32",x"33",x"34",x"35",x"36",x"37",x"38",x"39",x"3A",x"3B",x"3C",x"3D",x"3E",x"3F",
x"40",x"41",x"42",x"43",x"44",x"45",x"46",x"47",x"48",x"49",x"4A",x"4B",x"4C",x"4D",x"4E",x"4F",
x"50",x"51",x"52",x"53",x"54",x"55",x"56",x"57",x"58",x"59",x"5A",x"5B",x"5C",x"5D",x"5E",x"5F",
x"60",x"61",x"62",x"63",x"64",x"65",x"66",x"67",x"68",x"69",x"6A",x"6B",x"6C",x"6D",x"6E",x"6F",
x"70",x"71",x"72",x"73",x"74",x"75",x"76",x"77",x"78",x"79",x"7A",x"7B",x"7C",x"7D",x"7E",x"7F",
x"00",x"01",x"02",x"03",x"04",x"05",x"06",x"07",x"08",x"09",x"0A",x"0B",x"0C",x"0D",x"0E",x"0F",
x"10",x"11",x"12",x"13",x"14",x"15",x"16",x"17",x"18",x"19",x"1A",x"1B",x"1C",x"1D",x"1E",x"1F",
x"20",x"21",x"22",x"23",x"24",x"25",x"26",x"27",x"28",x"29",x"2A",x"2B",x"2C",x"2D",x"2E",x"2F",
x"30",x"31",x"32",x"33",x"34",x"35",x"36",x"37",x"38",x"39",x"3A",x"3B",x"3C",x"3D",x"3E",x"3F",
x"40",x"41",x"42",x"43",x"44",x"45",x"46",x"47",x"48",x"49",x"4A",x"4B",x"4C",x"4D",x"4E",x"4F",
x"50",x"51",x"52",x"53",x"54",x"55",x"56",x"57",x"58",x"59",x"5A",x"5B",x"5C",x"5D",x"5E",x"5F",
x"60",x"61",x"62",x"63",x"64",x"65",x"66",x"67",x"68",x"69",x"6A",x"6B",x"6C",x"6D",x"6E",x"6F",
x"70",x"71",x"72",x"73",x"74",x"75",x"76",x"77",x"78",x"79",x"7A",x"7B",x"7C",x"7D",x"7E",x"7F",

x"00",x"01",x"02",x"03",x"04",x"05",x"06",x"07",x"08",x"09",x"0A",x"0B",x"0C",x"0D",x"0E",x"0F",
x"10",x"11",x"12",x"13",x"14",x"15",x"16",x"17",x"18",x"19",x"1A",x"1B",x"1C",x"1D",x"1E",x"1F",
x"20",x"21",x"22",x"23",x"24",x"25",x"26",x"27",x"28",x"29",x"2A",x"2B",x"2C",x"2D",x"2E",x"2F",
x"30",x"31",x"32",x"33",x"34",x"35",x"36",x"37",x"38",x"39",x"3A",x"3B",x"3C",x"3D",x"3E",x"3F",
x"40",x"41",x"42",x"43",x"44",x"45",x"46",x"47",x"48",x"49",x"4A",x"4B",x"4C",x"4D",x"4E",x"4F",
x"50",x"51",x"52",x"53",x"54",x"55",x"56",x"57",x"58",x"59",x"5A",x"5B",x"5C",x"5D",x"5E",x"5F",
x"60",x"61",x"62",x"63",x"64",x"65",x"66",x"67",x"68",x"69",x"6A",x"6B",x"6C",x"6D",x"6E",x"6F",
x"70",x"71",x"72",x"73",x"74",x"75",x"76",x"77",x"78",x"79",x"7A",x"7B",x"7C",x"7D",x"7E",x"7F",
x"00",x"01",x"02",x"03",x"04",x"05",x"06",x"07",x"08",x"09",x"0A",x"0B",x"0C",x"0D",x"0E",x"0F",
x"10",x"11",x"12",x"13",x"14",x"15",x"16",x"17",x"18",x"19",x"1A",x"1B",x"1C",x"1D",x"1E",x"1F",
x"20",x"21",x"22",x"23",x"24",x"25",x"26",x"27",x"28",x"29",x"2A",x"2B",x"2C",x"2D",x"2E",x"2F",
x"30",x"31",x"32",x"33",x"34",x"35",x"36",x"37",x"38",x"39",x"3A",x"3B",x"3C",x"3D",x"3E",x"3F",
x"40",x"41",x"42",x"43",x"44",x"45",x"46",x"47",x"48",x"49",x"4A",x"4B",x"4C",x"4D",x"4E",x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"20",
x"20",
x"20",
x"20",
x"53",
x"55",
x"48",
x"41",
x"53",
x"48",
x"4B",
x"41",
x"20",
x"20",
x"20",
x"20",
x"53",
x"56",
x"49",
x"4E",
x"20",
x"20",
x"20",
x"20",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"20",
x"20",
x"20",
x"20",
x"53",
x"55",
x"48",
x"41",
x"53",
x"48",
x"4B",
x"41",
x"20",
x"20",
x"20",
x"20",
x"53",
x"56",
x"49",
x"4E",
x"20",
x"20",
x"20",
x"20",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"20",
x"20",
x"20",
x"20",
x"53",
x"55",
x"48",
x"41",
x"53",
x"48",
x"4B",
x"41",
x"20",
x"20",
x"20",
x"20",
x"53",
x"56",
x"49",
x"4E",
x"20",
x"20",
x"20",
x"20",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"20",
x"20",
x"20",
x"20",
x"53",
x"55",
x"48",
x"41",
x"53",
x"48",
x"4B",
x"41",
x"20",
x"20",
x"20",
x"20",
x"53",
x"56",
x"49",
x"4E",
x"20",
x"20",
x"20",
x"20",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F",
x"00",
x"01",
x"02",
x"03",
x"04",
x"05",
x"06",
x"07",
x"08",
x"09",
x"0A",
x"0B",
x"0C",
x"0D",
x"0E",
x"0F",
x"10",
x"11",
x"12",
x"13",
x"14",
x"15",
x"16",
x"17",
x"18",
x"19",
x"1A",
x"1B",
x"1C",
x"1D",
x"1E",
x"1F",
x"20",
x"21",
x"22",
x"23",
x"24",
x"25",
x"26",
x"27",
x"28",
x"29",
x"2A",
x"2B",
x"2C",
x"2D",
x"2E",
x"2F",
x"30",
x"31",
x"32",
x"33",
x"34",
x"35",
x"36",
x"37",
x"38",
x"39",
x"3A",
x"3B",
x"3C",
x"3D",
x"3E",
x"3F",
x"40",
x"41",
x"42",
x"43",
x"44",
x"45",
x"46",
x"47",
x"48",
x"49",
x"4A",
x"4B",
x"4C",
x"4D",
x"4E",
x"4F",
x"50",
x"51",
x"52",
x"53",
x"54",
x"55",
x"56",
x"57",
x"58",
x"59",
x"5A",
x"5B",
x"5C",
x"5D",
x"5E",
x"5F",
x"60",
x"61",
x"62",
x"63",
x"64",
x"65",
x"66",
x"67",
x"68",
x"69",
x"6A",
x"6B",
x"6C",
x"6D",
x"6E",
x"6F",
x"70",
x"71",
x"72",
x"73",
x"74",
x"75",
x"76",
x"77",
x"78",
x"79",
x"7A",
x"7B",
x"7C",
x"7D",
x"7E",
x"7F"
	);
--    attribute syn_romstyle : string;
--    attribute syn_romstyle of ROM: signal is "black_rom";


	signal RAM_SCREEN_Hi: ram_type := (   -- 2^13-by-16
x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",
x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",
x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",
x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",
x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",
x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",
x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",
x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",
x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",
x"14",x"14",x"14",x"14",x"14",x"14",x"14",x"14",x"14",x"14",x"14",x"14",x"14",x"14",x"14",x"14",
x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"15",
x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",
x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",
x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",

x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"63",
x"63",
x"63",
x"63",
x"63",
x"63",
x"63",
x"63",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"63",
x"63",
x"63",
x"63",
x"63",
x"63",
x"63",
x"63",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"63",
x"63",
x"63",
x"63",
x"63",
x"63",
x"63",
x"63",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"63",
x"63",
x"63",
x"63",
x"63",
x"63",
x"63",
x"63",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"10",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"12",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"13",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"14",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"15",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"16",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"17",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"1F",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"21",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"23",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"24",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"25",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"26",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"27",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"2F",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"31",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"32",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"34",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"35",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"36",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"37",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"3F",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"41",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"42",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"43",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"45",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"46",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"47",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"4F",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"51",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"52",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"53",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"54",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"55",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"56",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"57",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"5F",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"61",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"63",
x"63",
x"63",
x"63",
x"63",
x"63",
x"63",
x"63",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"64",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"65",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"66",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"67",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"6F",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"71",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"72",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"73",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"74",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"75",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"76",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"77",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"7F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"05",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"06",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"07",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F",
x"0F"
	);


--------------------------------------------------------------------------
-- FONT Table                                                           --
--------------------------------------------------------------------------

--------------------------------------------------------------------------
-- FONT lo byte                                                         --
--------------------------------------------------------------------------
	type rom_type is array (0 to 4095) of std_logic_vector(7 downto 0);
	signal RAM_FONT8_Lo: rom_type := (
--------------------------------------------------------------------------
-- FONT 8x8 1 bit on pixel (2048 bytes)                                --
--------------------------------------------------------------------------
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",

"00011100",
"00100010",
"01010101",
"01000001",
"01010101",
"01001001",
"00100010",
"00011100",

"00011100",
"00111110",
"01001001",
"01111111",
"01001001",
"01100011",
"00111110",
"00011100",

"00000000",
"00110110",
"01001001",
"01000001",
"00100010",
"00010100",
"00001000",
"00000000",

"00001000",
"00010100",
"00100010",
"01000001",
"00100010",
"00010100",
"00001000",
"00000000",

"00001000",
"00010100",
"00001000",
"00100010",
"01010101",
"00100010",
"00001000",
"00011100",

"00001000",
"00010100",
"00100010",
"01000001",
"01001001",
"00110110",
"00001000",
"00011100",

"00000000",
"00000000",
"00000000",
"00011100",
"00011100",
"00000000",
"00000000",
"00000000",

"01111111",
"01111111",
"01111111",
"01100011",
"01100011",
"01111111",
"01111111",
"01111111",

"00000000",
"00000000",
"00011100",
"00100010",
"00100010",
"00011100",
"00000000",
"00000000",

"01111111",
"01111111",
"01100011",
"01011101",
"01011101",
"01100011",
"01111111",
"01111111",

"00000000",
"00001110",
"00000110",
"00001010",
"00110000",
"01001000",
"00110000",
"00000000",

"00011100",
"00100010",
"00100010",
"00011100",
"00001000",
"00001000",
"00011100",
"00001000",

"00001100",
"00001110",
"00001010",
"00001010",
"00001000",
"00111000",
"00111000",
"00000000",

"00011111",
"00010001",
"00011111",
"00010001",
"00010111",
"01110111",
"01110000",
"00000000",

"00000000",
"00101010",
"00011100",
"00110110",
"00011100",
"00101010",
"00000000",
"00000000",

"00000000",
"00000000",
"00100000",
"00111000",
"00111110",
"00111000",
"00100000",
"00000000",

"00000000",
"00000000",
"00000010",
"00001110",
"00111110",
"00001110",
"00000010",
"00000000",

"00000000",
"00010000",
"00111000",
"00010000",
"00010000",
"00111000",
"00010000",
"00000000",

"00000000",
"00100100",
"00100100",
"00100100",
"00100100",
"00000000",
"00100100",
"00000000",

"00000000",
"01111110",
"10100100",
"01100100",
"00100100",
"00100100",
"00100100",
"00000000",

"00000000",
"00111100",
"01000000",
"00111100",
"01000010",
"00111100",
"00000010",
"00111100",

"00000000",
"00000000",
"00000000",
"11111110",
"11111110",
"00000000",
"00000000",
"00000000",

"00000000",
"00010000",
"00111000",
"00010000",
"00010000",
"00111000",
"00010000",
"01111100",

"00000000",
"00010000",
"00111000",
"00010000",
"00010000",
"00010000",
"00010000",
"00000000",

"00000000",
"00010000",
"00010000",
"00010000",
"00010000",
"00111000",
"00010000",
"00000000",

"00000000",
"00000000",
"00001000",
"00000100",
"01111110",
"00000100",
"00001000",
"00000000",

"00000000",
"00000000",
"00010000",
"00100000",
"01111110",
"00100000",
"00010000",
"00000000",

"00000000",
"00000000",
"01000000",
"01000000",
"01111110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"01000100",
"11111110",
"01000100",
"00000000",
"00000000",
"00000000",
"00000000",
"00010000",
"00111000",
"01111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"01111100",
"00111000",
"00010000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001000",
"00001000",
"00001000",
"00001000",
"00000000",
"00001000",
"00000000",
"00000000",
"00100100",
"00100100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00100100",
"01111110",
"00100100",
"01111110",
"00100100",
"00000000",
"00000000",
"00010000",
"01111100",
"10010000",
"01111100",
"00010010",
"01111100",
"00010000",
"00000000",
"01100010",
"01100100",
"00001000",
"00010000",
"00100110",
"01000110",
"00000000",
"00000000",
"00011000",
"00100100",
"00011000",
"00101010",
"01000100",
"00111010",
"00000000",
"00000000",
"00011000",
"00001000",
"00010000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001000",
"00010000",
"00010000",
"00010000",
"00010000",
"00001000",
"00000000",
"00000000",
"00010000",
"00001000",
"00001000",
"00001000",
"00001000",
"00010000",
"00000000",
"00000000",
"01000100",
"00101000",
"01111100",
"00101000",
"01000100",
"00000000",
"00000000",
"00000000",
"00010000",
"00010000",
"01111100",
"00010000",
"00010000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00011000",
"00001000",
"00010000",
"00000000",
"00000000",
"00000000",
"00000000",
"01111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00011000",
"00011000",
"00000000",
"00000000",
"00001000",
"00001000",
"00010000",
"00010000",
"00100000",
"00100000",
"00000000",
"00000000",

"00111100",
"01000110",
"01001010",
"01010010",
"01100010",
"00111100",
"00000000",
"00000000",

"00001000",
"00011000",
"00101000",
"00001000",
"00001000",
"00111110",
"00000000",
"00000000",
"00111100",
"01000010",
"00000010",
"00111100",
"01000000",
"01111110",
"00000000",
"00000000",
"01111110",
"00000100",
"00001000",
"00000100",
"01000010",
"00111100",
"00000000",
"00000000",
"00001000",
"00010000",
"00100100",
"01111110",
"00000100",
"00001110",
"00000000",
"00000000",
"01111110",
"01000000",
"01111100",
"00000010",
"01000010",
"00111100",
"00000000",
"00000000",
"00111100",
"01000000",
"01111100",
"01000010",
"01000010",
"00111100",
"00000000",
"00000000",
"01111110",
"01000010",
"00000100",
"00001000",
"00010000",
"00100000",
"00000000",
"00000000",
"00111100",
"01000010",
"00111100",
"01000010",
"01000010",
"00111100",
"00000000",
"00000000",
"00111100",
"01000010",
"01000010",
"00111110",
"00000010",
"00111100",
"00000000",
"00000000",
"00000000",
"00001100",
"00001100",
"00000000",
"00001100",
"00001100",
"00000000",
"00000000",
"00000000",
"00011000",
"00011000",
"00000000",
"00011000",
"00001000",
"00010000",
"00000000",
"00000000",
"00011000",
"00110000",
"01100000",
"00110000",
"00011000",
"00000000",
"00000000",
"00000000",
"00000000",
"01111110",
"00000000",
"01111110",
"00000000",
"00000000",
"00000000",
"00000000",
"00110000",
"00011000",
"00001100",
"00011000",
"00110000",
"00000000",
"00000000",
"00111000",
"01000100",
"00001000",
"00010000",
"00000000",
"00010000",
"00000000",

"00111100",
"01000010",
"10011110",
"10100010",
"10100010",
"10011110",
"01000000",
"00111100",

"00000000",
"00011000",
"00100100",
"01000010",
"01111110",
"01000010",
"11100110",
"00000000",
"00000000",
"01111100",
"00100010",
"00111100",
"00100010",
"00100010",
"01111100",
"00000000",
"00000000",
"00111110",
"01000010",
"01000000",
"01000000",
"01000010",
"00111100",
"00000000",
"00000000",
"01111100",
"00100010",
"00100010",
"00100010",
"00100010",
"01111100",
"00000000",
"00000000",
"01111110",
"00100000",
"00111100",
"00100000",
"00100000",
"01111110",
"00000000",
"00000000",
"01111110",
"00100000",
"00111100",
"00100000",
"00100000",
"01110000",
"00000000",
"00000000",
"00111100",
"01000010",
"01000000",
"01001110",
"01000010",
"00111100",
"00000000",
"00000000",
"11101110",
"01000100",
"01111100",
"01000100",
"01000100",
"11101110",
"00000000",
"00000000",
"01111100",
"00010000",
"00010000",
"00010000",
"00010000",
"01111100",
"00000000",
"00000000",
"00111110",
"00001000",
"00001000",
"00001000",
"01001000",
"00110000",
"00000000",
"00000000",
"11101110",
"01001000",
"01110000",
"01001000",
"01000100",
"11101110",
"00000000",
"00000000",
"01000000",
"01000000",
"01000000",
"01000000",
"01000100",
"01111100",
"00000000",
"00000000",
"11000110",
"11000110",
"10101010",
"10010010",
"10000010",
"11000110",
"00000000",
"00000000",
"01000010",
"01100010",
"01010010",
"01001010",
"01000110",
"11000010",
"00000000",
"00000000",
"00111100",
"01000010",
"01000010",
"01000010",
"01000010",
"00111100",
"00000000",
"00000000",
"11111000",
"01000100",
"01000100",
"01111000",
"01000000",
"11100000",
"00000000",
"00000000",
"00111100",
"01000010",
"01000010",
"01001010",
"01000100",
"00111010",
"00000000",
"00000000",
"11111000",
"01000100",
"01000100",
"01111000",
"01001000",
"11100110",
"00000000",
"00000000",
"00111100",
"01000000",
"00111100",
"00000010",
"01000010",
"00111100",
"00000000",
"00000000",
"11111110",
"10010010",
"00010000",
"00010000",
"00010000",
"00111000",
"00000000",
"00000000",
"11100110",
"01000010",
"01000010",
"01000010",
"01000010",
"00111100",
"00000000",
"00000000",
"11000110",
"10000010",
"01000100",
"01000100",
"00101000",
"00010000",
"00000000",
"00000000",
"11000110",
"10000010",
"10010010",
"10010010",
"01101100",
"01000100",
"00000000",
"00000000",
"11000110",
"00101000",
"00010000",
"00101000",
"01000100",
"11000110",
"00000000",
"00000000",
"11000110",
"01000100",
"00101000",
"00010000",
"00010000",
"00111000",
"00000000",
"00000000",
"01111110",
"01000100",
"00001000",
"00010000",
"00100010",
"01111110",
"00000000",
"00000000",
"00011100",
"00010000",
"00010000",
"00010000",
"00010000",
"00011100",
"00000000",
"00000000",
"00100000",
"00010000",
"00010000",
"00001000",
"00001000",
"00000100",
"00000000",
"00000000",
"00111000",
"00001000",
"00001000",
"00001000",
"00001000",
"00111000",
"00000000",
"00000000",
"00001000",
"00010100",
"00100010",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"00010000",
"00001000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111000",
"00000100",
"00111100",
"01000100",
"00111010",
"00000000",
"00000000",
"01100000",
"00100000",
"00111100",
"00100010",
"00100010",
"01111100",
"00000000",
"00000000",
"00000000",
"00111110",
"01000010",
"01000000",
"01000010",
"00111100",
"00000000",
"00000000",
"00000110",
"00000100",
"00111100",
"01000100",
"01000100",
"00111110",
"00000000",
"00000000",
"00000000",
"00111100",
"01000010",
"01111110",
"01000000",
"00111100",
"00000000",
"00000000",
"00001100",
"00010000",
"00111000",
"00010000",
"00010000",
"00111000",
"00000000",
"00000000",
"00000000",
"00111100",
"01000010",
"01000010",
"00111110",
"00000010",
"00111100",
"00000000",
"11000000",
"01000000",
"01111100",
"01000010",
"01000010",
"11100110",
"00000000",
"00000000",
"00001000",
"00000000",
"00011000",
"00001000",
"00001000",
"00011100",
"00000000",
"00000000",
"00001000",
"00000000",
"00011100",
"00001000",
"00001000",
"01001000",
"00110000",
"00000000",
"11000000",
"01000000",
"01000110",
"01111000",
"01000100",
"11100110",
"00000000",
"00000000",
"00110000",
"00010000",
"00010000",
"00010000",
"00010000",
"00111000",
"00000000",
"00000000",
"00000000",
"10101100",
"11010010",
"10010010",
"10010010",
"10010010",
"00000000",
"00000000",
"00000000",
"11011100",
"01100010",
"01000010",
"01000010",
"11100010",
"00000000",
"00000000",
"00000000",
"00111100",
"01000010",
"01000010",
"01000010",
"00111100",
"00000000",
"00000000",
"00000000",
"01111100",
"00100010",
"00100010",
"00111100",
"00100000",
"01110000",
"00000000",
"00000000",
"00111110",
"01000100",
"01000100",
"00111100",
"00000100",
"00000110",
"00000000",
"00000000",
"01101100",
"00110010",
"00100000",
"00100000",
"01110000",
"00000000",
"00000000",
"00000000",
"00111100",
"01000000",
"00111100",
"00000010",
"00111100",
"00000000",
"00000000",
"00010000",
"00010000",
"00111000",
"00010000",
"00010000",
"00001100",
"00000000",
"00000000",
"00000000",
"11001110",
"01000100",
"01000100",
"01000100",
"00111010",
"00000000",
"00000000",
"00000000",
"11101110",
"01000100",
"00101000",
"00101000",
"00010000",
"00000000",
"00000000",
"00000000",
"11000110",
"10000010",
"10010010",
"10101010",
"01000100",
"00000000",
"00000000",
"00000000",
"11100110",
"00100100",
"00011000",
"00100100",
"11100110",
"00000000",
"00000000",
"00000000",
"11000110",
"00100100",
"00100100",
"00011000",
"00010000",
"01100000",
"00000000",
"00000000",
"01111110",
"00000100",
"00011000",
"00100000",
"01111110",
"00000000",
"00000000",
"00001000",
"00010000",
"00010000",
"00110000",
"00010000",
"00010000",
"00001000",
"00000000",
"00001000",
"00001000",
"00001000",
"00000000",
"00001000",
"00001000",
"00001000",
"00000000",
"00010000",
"00001000",
"00001000",
"00001100",
"00001000",
"00001000",
"00010000",
"00000000",
"00000000",
"00110000",
"01001001",
"00000110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00010000",
"00101000",
"01111100",
"00000000",
"00000000",
"00111000",
"01000100",
"01000100",
"01111100",
"01000100",
"11001110",
"00000000",
"00000000",
"01111100",
"00100000",
"00111100",
"00100010",
"00100010",
"01111100",
"00000000",
"00000000",
"01111100",
"00100010",
"00111100",
"00100010",
"00100010",
"01111100",
"00000000",
"00000000",
"00111110",
"00010010",
"00010000",
"00010000",
"00010000",
"00111000",
"00000000",
"00000000",
"00011110",
"00100100",
"00100100",
"00100100",
"00100100",
"01111110",
"01000010",
"00000000",
"01111110",
"00100010",
"00111000",
"00100000",
"00100010",
"01111110",
"00000000",
"00000000",
"11010110",
"01010100",
"00111000",
"01010100",
"10010010",
"10010010",
"00000000",
"00000000",
"00111100",
"01000010",
"00001100",
"00000010",
"01000010",
"00111100",
"00000000",
"00000000",
"01000010",
"01000110",
"01001010",
"01010010",
"01100010",
"01000010",
"00000000",
"00011000",
"01000010",
"01000110",
"01001010",
"01010010",
"01100010",
"01000010",
"00000000",
"00000000",
"01100100",
"00101000",
"00110000",
"00101000",
"00100100",
"01100110",
"00000000",
"00000000",
"00001110",
"00010010",
"00100010",
"00100010",
"00100010",
"01100010",
"00000000",
"00000000",
"11000110",
"01101100",
"01010100",
"01010100",
"01000100",
"11101110",
"00000000",
"00000000",
"11101110",
"01000100",
"01111100",
"01000100",
"01000100",
"11101110",
"00000000",
"00000000",
"00111100",
"01000010",
"01000010",
"01000010",
"01000010",
"00111100",
"00000000",
"00000000",
"11111110",
"01000100",
"01000100",
"01000100",
"01000100",
"11101110",
"00000000",
"00000000",
"01111100",
"00100010",
"00100010",
"00111100",
"00100000",
"01110000",
"00000000",
"00000000",
"00111100",
"01000010",
"01000000",
"01000000",
"01000010",
"00111100",
"00000000",
"00000000",
"01111100",
"01010100",
"00010000",
"00010000",
"00010000",
"00111000",
"00000000",
"00000000",
"11000110",
"01000100",
"00100100",
"00011000",
"00001000",
"01110000",
"00000000",
"00000000",
"00010000",
"01111100",
"10010010",
"10010010",
"10010010",
"01111100",
"00010000",
"00000000",
"01100110",
"00100100",
"00011000",
"00011000",
"00100100",
"01100110",
"00000000",
"00000000",
"11101110",
"01000100",
"01000100",
"01000100",
"01000100",
"11111110",
"00000010",
"00000000",
"11101110",
"01000100",
"01000100",
"00111100",
"00000100",
"00001110",
"00000000",
"00000000",
"10010010",
"10010010",
"10010010",
"10010010",
"10010010",
"11111110",
"00000000",
"00000000",
"10010010",
"10010010",
"10010010",
"10010010",
"10010010",
"11111111",
"00000001",
"00000000",
"11100000",
"10100000",
"00111100",
"00100010",
"00100010",
"01111100",
"00000000",
"00000000",
"11100010",
"01000010",
"01110010",
"01001010",
"01001010",
"11110010",
"00000000",
"00000000",
"01110000",
"00100000",
"00111100",
"00100010",
"00100010",
"01111100",
"00000000",
"00000000",
"00111100",
"01000010",
"00011110",
"00000010",
"01000010",
"00111100",
"00000000",
"00000000",
"10011100",
"10100010",
"10100010",
"11100010",
"10100010",
"10011100",
"00000000",
"00000000",
"00111110",
"01000100",
"01000100",
"00111100",
"00010100",
"01100110",
"00000000",
"00000000",
"00000000",
"00111000",
"00000100",
"00111100",
"01000100",
"00111010",
"00000000",
"00000010",
"00111100",
"01000000",
"00111100",
"01000010",
"01000010",
"00111100",
"00000000",
"00000000",
"00000000",
"01111100",
"00100010",
"00111100",
"00100010",
"01111100",
"00000000",
"00000000",
"00000000",
"01111110",
"00100010",
"00100000",
"00100000",
"01110000",
"00000000",
"00000000",
"00000000",
"00111110",
"00010100",
"00100100",
"00100100",
"01111110",
"01000010",
"00000000",
"00000000",
"00111100",
"01000010",
"01111110",
"01000000",
"00111100",
"00000000",
"00000000",
"00000000",
"11010110",
"01010100",
"00111000",
"01010100",
"11010110",
"00000000",
"00000000",
"00000000",
"00111100",
"01000010",
"00001100",
"01000010",
"00111100",
"00000000",
"00000000",
"00000000",
"11100110",
"01000110",
"01001010",
"01010010",
"11100110",
"00000000",
"00011000",
"00000000",
"11100110",
"01000110",
"01001010",
"01010010",
"11100110",
"00000000",
"00000000",
"00000000",
"11100110",
"01001000",
"01110000",
"01001000",
"11100110",
"00000000",
"00000000",
"00000000",
"00111110",
"00010100",
"00010100",
"00100100",
"01101110",
"00000000",
"00000000",
"00000000",
"11000110",
"11000110",
"10101010",
"10010010",
"10000010",
"00000000",
"00000000",
"00000000",
"11101110",
"01000100",
"01111100",
"01000100",
"11101110",
"00000000",
"00000000",
"00000000",
"00111100",
"01000010",
"01000010",
"01000010",
"00111100",
"00000000",
"00000000",
"00000000",
"11111110",
"01000100",
"01000100",
"01000100",
"11101110",
"00000000",
"10001000",
"00100010",
"10001000",
"00100010",
"10001000",
"00100010",
"10001000",
"00100010",
"10010010",
"01001001",
"10010010",
"01001001",
"10010010",
"01001001",
"10010010",
"00000000",
"10101010",
"01010101",
"10101010",
"01010101",
"10101010",
"01010101",
"10101010",
"00000000",
"00010000",
"00010000",
"00010000",
"00010000",
"00010000",
"00010000",
"00010000",
"00010000",
"00010000",
"00010000",
"00010000",
"11110000",
"00010000",
"00010000",
"00010000",
"00010000",
"00010000",
"00010000",
"11110000",
"00010000",
"11110000",
"00010000",
"00010000",
"00010000",
"00101000",
"00101000",
"00101000",
"11101000",
"00101000",
"00101000",
"00101000",
"00101000",
"00000000",
"00000000",
"00000000",
"11111000",
"00101000",
"00101000",
"00101000",
"00101000",
"00000000",
"00000000",
"11110000",
"00010000",
"11110000",
"00010000",
"00010000",
"00010000",
"00101000",
"00101000",
"11101000",
"00001000",
"11101000",
"00101000",
"00101000",
"00101000",
"00101000",
"00101000",
"00101000",
"00101000",
"00101000",
"00101000",
"00101000",
"00101000",
"00000000",
"00000000",
"11111000",
"00001000",
"11101000",
"00101000",
"00101000",
"00101000",
"00101000",
"00101000",
"11101000",
"00001000",
"11111000",
"00000000",
"00000000",
"00000000",
"00101000",
"00101000",
"00101000",
"11111000",
"00000000",
"00000000",
"00000000",
"00000000",
"00010000",
"00010000",
"11110000",
"00010000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00010000",
"00010000",
"00010000",
"00010000",
"00010000",
"00010000",
"00010000",
"00011111",
"00000000",
"00000000",
"00000000",
"00000000",
"00010000",
"00010000",
"00010000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00010000",
"00010000",
"00010000",
"00010000",
"00010000",
"00010000",
"00010000",
"00011111",
"00010000",
"00010000",
"00010000",
"00010000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00010000",
"00010000",
"00010000",
"11111111",
"00010000",
"00010000",
"00010000",
"00010000",
"00010000",
"00010000",
"00011111",
"00010000",
"00011111",
"00010000",
"00010000",
"00010000",
"00101000",
"00101000",
"00101000",
"00101111",
"00101000",
"00101000",
"00101000",
"00101000",
"00101000",
"00101000",
"00101111",
"00100000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"00100000",
"00101111",
"00101000",
"00101000",
"00101000",
"00101000",
"00101000",
"11101111",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"11101111",
"00101000",
"00101000",
"00101000",
"00101000",
"00101000",
"00101111",
"00100000",
"00101111",
"00101000",
"00101000",
"00101000",
"00000000",
"00000000",
"11111111",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00101000",
"00101000",
"11101111",
"00000000",
"11101111",
"00101000",
"00101000",
"00101000",
"00010000",
"00010000",
"11111111",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00101000",
"00101000",
"00101000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"11111111",
"00010000",
"00010000",
"00010000",
"00000000",
"00000000",
"00000000",
"11111111",
"00101000",
"00101000",
"00101000",
"00101000",
"00101000",
"00101000",
"00101000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00010000",
"00010000",
"00011111",
"00010000",
"00011111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00011111",
"00010000",
"00011111",
"00010000",
"00010000",
"00010000",
"00000000",
"00000000",
"00000000",
"00111111",
"00101000",
"00101000",
"00101000",
"00101000",
"00101000",
"00101000",
"00101000",
"11101111",
"00101000",
"00101000",
"00101000",
"00101000",
"00010000",
"00010000",
"11111111",
"00000000",
"11111111",
"00010000",
"00010000",
"00010000",
"00010000",
"00010000",
"00010000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00011111",
"00010000",
"00010000",
"00010000",
"00010000",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"11111111",
"11111111",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"11111111",
"11111111",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"01111100",
"00100010",
"00100010",
"00111100",
"00100000",
"01110000",
"00000000",
"00000000",
"00111100",
"01000010",
"01000000",
"01000010",
"00111100",
"00000000",
"00000000",
"00000000",
"01111100",
"01010100",
"00010000",
"00010000",
"00111000",
"00000000",
"00000000",
"00000000",
"11101110",
"01000100",
"01000100",
"00111100",
"00000100",
"01111000",
"00000000",
"00000000",
"00010000",
"01111100",
"10010010",
"10010010",
"01111100",
"00010000",
"00000000",
"00000000",
"11100110",
"00100100",
"00011000",
"00100100",
"11100110",
"00000000",
"00000000",
"00000000",
"11101110",
"01000100",
"01000100",
"01000100",
"11111110",
"00000010",
"00000000",
"00000000",
"11101110",
"01000100",
"00111100",
"00000100",
"00001110",
"00000000",
"00000000",
"00000000",
"10010010",
"10010010",
"10010010",
"10010010",
"11111110",
"00000000",
"00000000",
"00000000",
"10010010",
"10010010",
"10010010",
"10010010",
"11111110",
"00000010",
"00000000",
"00000000",
"11100000",
"10100000",
"00111100",
"00100010",
"01111100",
"00000000",
"00000000",
"00000000",
"11100010",
"01000010",
"01110010",
"01001010",
"11110010",
"00000000",
"00000000",
"00000000",
"01110000",
"00100000",
"00111100",
"00100010",
"01111100",
"00000000",
"00000000",
"00000000",
"00111100",
"01000010",
"00011110",
"01000010",
"00111100",
"00000000",
"00000000",
"00000000",
"10011100",
"10100010",
"11100010",
"10100010",
"10011100",
"00000000",
"00000000",
"00000000",
"00111110",
"01000100",
"00111100",
"00100100",
"01101110",
"00000000",
"00100100",
"01111110",
"00100010",
"00111000",
"00100000",
"00100010",
"01111110",
"00000000",
"00100100",
"00000000",
"00111100",
"01000010",
"01111110",
"01000000",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000110",
"00001100",
"00011000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"01100000",
"00110000",
"00011000",
"00011000",
"00110000",
"01100000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00011000",
"00001100",
"00000110",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001000",
"00000100",
"01111110",
"00000100",
"00001000",
"00000000",
"00000000",
"00000000",
"00010000",
"00100000",
"01111110",
"00100000",
"00010000",
"00000000",
"00000000",
"00010000",
"00111000",
"01010100",
"00010000",
"00010000",
"00010000",
"00000000",
"00000000",
"00010000",
"00010000",
"00010000",
"01010100",
"00111000",
"00010000",
"00000000",
"00000000",
"00011000",
"00000000",
"01111110",
"00000000",
"00011000",
"00000000",
"00000000",
"00010000",
"00010000",
"01111100",
"00010000",
"00010000",
"00000000",
"01111100",
"00000000",
"00000000",
"10001011",
"10001011",
"11001000",
"10101011",
"10011000",
"10001000",
"00000000",
"00000000",
"00000000",
"01000010",
"00111100",
"01000010",
"00111100",
"01000010",
"00000000",
"00000000",
"00000000",
"00000000",
"00011100",
"00011100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",

--------------------------------------------------------------
-- FONT 8x8 2 bits on pixel (2048 bytes)
--------------------------------------------------------------
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"00110011",
"00000011",
"00110011",
"11000011",
"00001100",
"11110000",
"11110000",
"11111100",
"11000011",
"11111111",
"11000011",
"00001111",
"11111100",
"11110000",
"00000000",
"00111100",
"11000011",
"00000011",
"00001100",
"00110000",
"11000000",
"00000000",
"11000000",
"00110000",
"00001100",
"00000011",
"00001100",
"00110000",
"11000000",
"00000000",
"11000000",
"00110000",
"11000000",
"00001100",
"00110011",
"00001100",
"11000000",
"11110000",
"11000000",
"00110000",
"00001100",
"00000011",
"11000011",
"00111100",
"11000000",
"11110000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"11111111",
"00001111",
"00001111",
"11111111",
"11111111",
"11111111",
"00000000",
"00000000",
"11110000",
"00001100",
"00001100",
"11110000",
"00000000",
"00000000",
"11111111",
"11111111",
"00001111",
"11110011",
"11110011",
"00001111",
"11111111",
"11111111",
"00000000",
"11111100",
"00111100",
"11001100",
"00000000",
"11000000",
"00000000",
"00000000",
"11110000",
"00001100",
"00001100",
"11110000",
"11000000",
"11000000",
"11110000",
"11000000",
"11110000",
"11111100",
"11001100",
"11001100",
"11000000",
"11000000",
"11000000",
"00000000",
"11111111",
"00000011",
"11111111",
"00000011",
"00111111",
"00111111",
"00000000",
"00000000",
"00000000",
"11001100",
"11110000",
"00111100",
"11110000",
"11001100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11111100",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001100",
"11111100",
"11111100",
"11111100",
"00001100",
"00000000",
"00000000",
"00000000",
"11000000",
"00000000",
"00000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00110000",
"00110000",
"00110000",
"00110000",
"00000000",
"00110000",
"00000000",
"00000000",
"11111100",
"00110000",
"00110000",
"00110000",
"00110000",
"00110000",
"00000000",
"00000000",
"11110000",
"00000000",
"11110000",
"00001100",
"11110000",
"00001100",
"11110000",
"00000000",
"00000000",
"00000000",
"11111100",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"00000000",
"00000000",
"11000000",
"00000000",
"11110000",
"00000000",
"00000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"00110000",
"11111100",
"00110000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110000",
"11111100",
"00110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11000000",
"11000000",
"00000000",
"11000000",
"00000000",
"00000000",
"00110000",
"00110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110000",
"11111100",
"00110000",
"11111100",
"00110000",
"00000000",
"00000000",
"00000000",
"11110000",
"00000000",
"11110000",
"00001100",
"11110000",
"00000000",
"00000000",
"00001100",
"00110000",
"11000000",
"00000000",
"00111100",
"00111100",
"00000000",
"00000000",
"11000000",
"00110000",
"11000000",
"11001100",
"00110000",
"11001100",
"00000000",
"00000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00110000",
"11000000",
"11110000",
"11000000",
"00110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"00000000",
"00000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"11001100",
"00001100",
"00001100",
"11110000",
"00000000",
"00000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11111100",
"00000000",
"00000000",
"11110000",
"00001100",
"00001100",
"11110000",
"00000000",
"11111100",
"00000000",
"00000000",
"11111100",
"00110000",
"11000000",
"00110000",
"00001100",
"11110000",
"00000000",
"00000000",
"11000000",
"00000000",
"00110000",
"11111100",
"00110000",
"11111100",
"00000000",
"00000000",
"11111100",
"00000000",
"11110000",
"00001100",
"00001100",
"11110000",
"00000000",
"00000000",
"11110000",
"00000000",
"11110000",
"00001100",
"00001100",
"11110000",
"00000000",
"00000000",
"11111100",
"00001100",
"00110000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"11110000",
"00001100",
"00001100",
"11110000",
"00000000",
"00000000",
"11110000",
"00001100",
"00001100",
"11111100",
"00001100",
"11110000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"00000000",
"11110000",
"11110000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"00000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"11000000",
"00000000",
"00000000",
"00000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00000000",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11110000",
"11000000",
"00000000",
"00000000",
"00000000",
"11000000",
"00110000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"11111100",
"00001100",
"00001100",
"11111100",
"00000000",
"11110000",
"00000000",
"11000000",
"00110000",
"00001100",
"11111100",
"00001100",
"00111100",
"00000000",
"00000000",
"11110000",
"00001100",
"11110000",
"00001100",
"00001100",
"11110000",
"00000000",
"00000000",
"11111100",
"00001100",
"00000000",
"00000000",
"00001100",
"11110000",
"00000000",
"00000000",
"11110000",
"00001100",
"00001100",
"00001100",
"00001100",
"11110000",
"00000000",
"00000000",
"11111100",
"00000000",
"11110000",
"00000000",
"00000000",
"11111100",
"00000000",
"00000000",
"11111100",
"00000000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"00000000",
"11111100",
"00001100",
"11110000",
"00000000",
"00000000",
"11111100",
"00110000",
"11110000",
"00110000",
"00110000",
"11111100",
"00000000",
"00000000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00000000",
"00000000",
"11111100",
"11000000",
"11000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"11111100",
"11000000",
"00000000",
"11000000",
"00110000",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110000",
"11110000",
"00000000",
"00000000",
"00111100",
"00111100",
"11001100",
"00001100",
"00001100",
"00111100",
"00000000",
"00000000",
"00001100",
"00001100",
"00001100",
"11001100",
"00111100",
"00001100",
"00000000",
"00000000",
"11110000",
"00001100",
"00001100",
"00001100",
"00001100",
"11110000",
"00000000",
"00000000",
"11000000",
"00110000",
"00110000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"00001100",
"11001100",
"00110000",
"11001100",
"00000000",
"00000000",
"11000000",
"00110000",
"00110000",
"11000000",
"11000000",
"00111100",
"00000000",
"00000000",
"11110000",
"00000000",
"11110000",
"00001100",
"00001100",
"11110000",
"00000000",
"00000000",
"11111100",
"00001100",
"00000000",
"00000000",
"00000000",
"11000000",
"00000000",
"00000000",
"00111100",
"00001100",
"00001100",
"00001100",
"00001100",
"11110000",
"00000000",
"00000000",
"00111100",
"00001100",
"00110000",
"00110000",
"11000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00001100",
"00001100",
"00001100",
"11110000",
"00110000",
"00000000",
"00000000",
"00111100",
"11000000",
"00000000",
"11000000",
"00110000",
"00111100",
"00000000",
"00000000",
"00111100",
"00110000",
"11000000",
"00000000",
"00000000",
"11000000",
"00000000",
"00000000",
"11111100",
"00110000",
"11000000",
"00000000",
"00001100",
"11111100",
"00000000",
"00000000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"00110000",
"00000000",
"00000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"00000000",
"00000000",
"11000000",
"00110000",
"00001100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"00000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"00110000",
"11110000",
"00110000",
"11001100",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"00001100",
"11110000",
"00000000",
"00000000",
"00000000",
"11111100",
"00001100",
"00000000",
"00001100",
"11110000",
"00000000",
"00000000",
"00111100",
"00110000",
"11110000",
"00110000",
"00110000",
"11111100",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"11111100",
"00000000",
"11110000",
"00000000",
"00000000",
"11110000",
"00000000",
"11000000",
"00000000",
"00000000",
"11000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"00001100",
"11111100",
"00001100",
"11110000",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"00001100",
"00111100",
"00000000",
"00000000",
"11000000",
"00000000",
"11000000",
"11000000",
"11000000",
"11110000",
"00000000",
"00000000",
"11000000",
"00000000",
"11110000",
"11000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"11000000",
"00110000",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"00001100",
"00001100",
"00001100",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"00001100",
"00001100",
"00001100",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"00001100",
"00001100",
"11110000",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"00001100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00110000",
"00110000",
"11110000",
"00110000",
"00111100",
"00000000",
"00000000",
"11110000",
"00001100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00000000",
"11110000",
"00001100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"00000000",
"00000000",
"11110000",
"00000000",
"00000000",
"00000000",
"11111100",
"00110000",
"00110000",
"00110000",
"11001100",
"00000000",
"00000000",
"00000000",
"11111100",
"00110000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00001100",
"00001100",
"11001100",
"00110000",
"00000000",
"00000000",
"00000000",
"00111100",
"00110000",
"11000000",
"00110000",
"00111100",
"00000000",
"00000000",
"00000000",
"00111100",
"00110000",
"00110000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00110000",
"11000000",
"00000000",
"11111100",
"00000000",
"00000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"00000000",
"11000000",
"11000000",
"11000000",
"00000000",
"11000000",
"11000000",
"11000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11110000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000011",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11110000",
"00000000",
"00000000",
"11000000",
"00110000",
"00110000",
"11110000",
"00110000",
"11111100",
"00000000",
"00000000",
"11110000",
"00000000",
"11110000",
"00001100",
"00001100",
"11110000",
"00000000",
"00000000",
"11110000",
"00001100",
"11110000",
"00001100",
"00001100",
"11110000",
"00000000",
"00000000",
"11111100",
"00001100",
"00000000",
"00000000",
"00000000",
"11000000",
"00000000",
"00000000",
"11111100",
"00110000",
"00110000",
"00110000",
"00110000",
"11111100",
"00001100",
"00000000",
"11111100",
"00001100",
"11000000",
"00000000",
"00001100",
"11111100",
"00000000",
"00000000",
"00111100",
"00110000",
"11000000",
"00110000",
"00001100",
"00001100",
"00000000",
"00000000",
"11110000",
"00001100",
"11110000",
"00001100",
"00001100",
"11110000",
"00000000",
"00000000",
"00001100",
"00111100",
"11001100",
"00001100",
"00001100",
"00001100",
"00000000",
"11000000",
"00001100",
"00111100",
"11001100",
"00001100",
"00001100",
"00001100",
"00000000",
"00000000",
"00110000",
"11000000",
"00000000",
"11000000",
"00110000",
"00111100",
"00000000",
"00000000",
"11111100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00000000",
"00000000",
"00111100",
"11110000",
"00110000",
"00110000",
"00110000",
"11111100",
"00000000",
"00000000",
"11111100",
"00110000",
"11110000",
"00110000",
"00110000",
"11111100",
"00000000",
"00000000",
"11110000",
"00001100",
"00001100",
"00001100",
"00001100",
"11110000",
"00000000",
"00000000",
"11111100",
"00110000",
"00110000",
"00110000",
"00110000",
"11111100",
"00000000",
"00000000",
"11110000",
"00001100",
"00001100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"00000000",
"00000000",
"00001100",
"11110000",
"00000000",
"00000000",
"11110000",
"00110000",
"00000000",
"00000000",
"00000000",
"11000000",
"00000000",
"00000000",
"00111100",
"00110000",
"00110000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"00001100",
"00001100",
"11110000",
"00000000",
"00000000",
"00111100",
"00110000",
"11000000",
"11000000",
"00110000",
"00111100",
"00000000",
"00000000",
"11111100",
"00110000",
"00110000",
"00110000",
"00110000",
"11111100",
"00001100",
"00000000",
"11111100",
"00110000",
"00110000",
"11110000",
"00110000",
"11111100",
"00000000",
"00000000",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"11111100",
"00000000",
"00000000",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"11111111",
"00000011",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"00001100",
"11110000",
"00000000",
"00000000",
"00001100",
"00001100",
"00001100",
"11001100",
"11001100",
"00001100",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"00001100",
"11110000",
"00000000",
"00000000",
"11110000",
"00001100",
"11111100",
"00001100",
"00001100",
"11110000",
"00000000",
"00000000",
"11110000",
"00001100",
"00001100",
"00001100",
"00001100",
"11110000",
"00000000",
"00000000",
"11111100",
"00110000",
"00110000",
"11110000",
"00110000",
"00111100",
"00000000",
"00000000",
"00000000",
"11000000",
"00110000",
"11110000",
"00110000",
"11001100",
"00000000",
"00001100",
"11110000",
"00000000",
"11110000",
"00001100",
"00001100",
"11110000",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"11110000",
"00001100",
"11110000",
"00000000",
"00000000",
"00000000",
"11111100",
"00001100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00110000",
"00110000",
"00110000",
"11111100",
"00001100",
"00000000",
"00000000",
"11110000",
"00001100",
"11111100",
"00000000",
"11110000",
"00000000",
"00000000",
"00000000",
"00111100",
"00110000",
"11000000",
"00110000",
"00111100",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"11110000",
"00001100",
"11110000",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"11001100",
"00001100",
"00111100",
"00000000",
"11000000",
"00000000",
"00111100",
"00111100",
"11001100",
"00001100",
"00111100",
"00000000",
"00000000",
"00000000",
"00111100",
"11000000",
"00000000",
"11000000",
"00111100",
"00000000",
"00000000",
"00000000",
"11111100",
"00110000",
"00110000",
"00110000",
"11111100",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"11001100",
"00001100",
"00001100",
"00000000",
"00000000",
"00000000",
"11111100",
"00110000",
"11110000",
"00110000",
"11111100",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"00001100",
"00001100",
"11110000",
"00000000",
"00000000",
"00000000",
"11111100",
"00110000",
"00110000",
"00110000",
"11111100",
"00000000",
"11000000",
"00001100",
"11000000",
"00001100",
"11000000",
"00001100",
"11000000",
"00001100",
"00001100",
"11000011",
"00001100",
"11000011",
"00001100",
"11000011",
"00001100",
"00000000",
"11001100",
"00110011",
"11001100",
"00110011",
"11001100",
"00110011",
"11001100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11000000",
"11111111",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11111111",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"11111111",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11111111",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"11111111",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11111111",
"00000000",
"11111111",
"11000000",
"11000000",
"11000000",
"00000000",
"00000000",
"11111111",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11111111",
"00000000",
"11111111",
"11000000",
"11000000",
"11000000",
"00000000",
"00000000",
"11111111",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11111111",
"11000000",
"11000000",
"11000000",
"11000000",
"00000000",
"00000000",
"11111111",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"00001100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"00000000",
"00001100",
"11110000",
"00000000",
"00000000",
"00000000",
"11110000",
"00110000",
"00000000",
"00000000",
"11000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00110000",
"00110000",
"11110000",
"00110000",
"11000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"00001100",
"11110000",
"00000000",
"00000000",
"00000000",
"00111100",
"00110000",
"11000000",
"00110000",
"00111100",
"00000000",
"00000000",
"00000000",
"11111100",
"00110000",
"00110000",
"00110000",
"11111100",
"00001100",
"00000000",
"00000000",
"11111100",
"00110000",
"11110000",
"00110000",
"11111100",
"00000000",
"00000000",
"00000000",
"00001100",
"00001100",
"00001100",
"00001100",
"11111100",
"00000000",
"00000000",
"00000000",
"00001100",
"00001100",
"00001100",
"00001100",
"11111100",
"00001100",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"11110000",
"00000000",
"00000000",
"00000000",
"00001100",
"00001100",
"00001100",
"11001100",
"00001100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"11110000",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"11111100",
"00001100",
"11110000",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"00001100",
"00001100",
"11110000",
"00000000",
"00000000",
"00000000",
"11111100",
"00110000",
"11110000",
"00110000",
"11111100",
"00000000",
"00110000",
"11111100",
"00001100",
"11000000",
"00000000",
"00001100",
"11111100",
"00000000",
"00110000",
"00000000",
"11110000",
"00001100",
"11111100",
"00000000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00111100",
"11110000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11110000",
"00111100",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"00110000",
"11111100",
"00110000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"00110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110000",
"11000000",
"00000000",
"00000000",
"00000000",
"11000000",
"00000000",
"11111100",
"00000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00000000",
"00000000",
"00000000",
"11110000",
"00000000",
"00000000",
"11001111",
"11001111",
"11000000",
"11001111",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00001100",
"11110000",
"00001100",
"11110000",
"00001100",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000"
);

--------------------------------------------------------------
--
--------------------------------------------------------------
	signal RAM_FONT16_Lo: rom_type := (
--------------------------------------------------------------
---- FONT 16x16 1 bit on pixel or 8x16 2 bits on pixel (4096 bytes)
--------------------------------------------------------------
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00000011",
"00110011",
"00000011",
"00000011",
"11110011",
"11000011",
"00000011",
"00000011",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"11111111",
"11001111",
"11111111",
"11111111",
"00001111",
"00111111",
"11111111",
"11111111",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110000",
"11000000",
"00000000",
"00111100",
"11000011",
"00001100",
"00110000",
"11000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110000",
"11000000",
"00000000",
"00110011",
"00110011",
"00110011",
"00111111",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11110000",
"11110000",
"11000000",
"00111100",
"11111111",
"11111111",
"00111100",
"11000000",
"11110000",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11110000",
"11110000",
"11111100",
"11111111",
"11111111",
"11111111",
"11111100",
"11000000",
"11110000",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11110000",
"11110000",
"11110000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"11111111",
"11111111",
"00111111",
"00001111",
"00001111",
"00001111",
"00111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00001100",
"00001100",
"00001100",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"11111111",
"00001111",
"11000011",
"11110011",
"11110011",
"11110011",
"11000011",
"00001111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"00000000",
"11111100",
"11111100",
"11001100",
"00001100",
"11000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00111100",
"00111100",
"00111100",
"11110000",
"11000000",
"11111100",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00001111",
"00001111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00001111",
"00001111",
"11111111",
"00001111",
"00001111",
"00001111",
"00111111",
"00111111",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11001111",
"11110000",
"00111111",
"00111111",
"11110000",
"11001111",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11111100",
"11111100",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001100",
"00111100",
"11111100",
"11111100",
"11111100",
"11111100",
"11111100",
"11111100",
"00111100",
"00001100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11110000",
"11111100",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11111100",
"11110000",
"11000000",
"00000000",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00000000",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11001111",
"11001111",
"11001111",
"11001111",
"11001111",
"11001111",
"11001111",
"11001111",
"11001111",
"11001111",
"11001111",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00000000",
"11000000",
"11110000",
"00111100",
"00111100",
"11110000",
"11000000",
"11110000",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"11111100",
"11111100",
"11111100",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11110000",
"11111100",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11111100",
"11110000",
"11000000",
"11111100",
"00000000",
"00000000",
"00000000",
"11000000",
"11110000",
"11111100",
"11111111",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11111111",
"11111100",
"11110000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11110000",
"11111100",
"11111111",
"11111100",
"11110000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110000",
"00111100",
"11111111",
"00111100",
"00110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11110000",
"11110000",
"11111100",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"11111100",
"11110000",
"11110000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11110000",
"11111100",
"11111100",
"11111100",
"11111100",
"11110000",
"11000000",
"11000000",
"00000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00001111",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11111100",
"11111100",
"11110000",
"11110000",
"11110000",
"11111100",
"11111100",
"11110000",
"11110000",
"11110000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11111100",
"11001111",
"11001111",
"11000000",
"11000000",
"11111100",
"11001111",
"11001111",
"11001111",
"11001111",
"11111100",
"11000000",
"11000000",
"00000000",
"00000000",
"00111100",
"00111100",
"11110000",
"11110000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"11111100",
"11001100",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11110000",
"11110000",
"11110000",
"11000000",
"00111100",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11110000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"11110000",
"11111111",
"11111111",
"11110000",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11111100",
"11111100",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"11110000",
"11110000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00111100",
"11111100",
"11111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"10000000",
"10000000",
"10000000",
"10000000",
"10000000",
"10000000",
"10000000",
"10000000",
"10000000",
"10000000",
"10000000",
"10101000",
"00000000",
"00000000",
"00000000",
"00000000",
"01010000",
"00010100",
"00000101",
"00000101",
"00000101",
"00010100",
"01010000",
"01000000",
"00000000",
"00000000",
"00000101",
"01010101",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00111100",
"11110000",
"11000000",
"11110000",
"00111100",
"00001111",
"00001111",
"00001111",
"00001111",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110011",
"11111111",
"11110011",
"11110000",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00001111",
"00001111",
"00001111",
"00001111",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00111100",
"00000000",
"11110000",
"00111100",
"00001111",
"00001111",
"00001111",
"00001111",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00111100",
"00111100",
"11110000",
"11110000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00001111",
"00001111",
"00111100",
"11110000",
"00111100",
"00001111",
"00001111",
"00001111",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00001111",
"00001111",
"00001111",
"00001111",
"00111111",
"11111111",
"00001111",
"00001111",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00111100",
"11110000",
"11000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11110000",
"00111100",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"11111100",
"00000000",
"11111100",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11110000",
"00111100",
"11110000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00001111",
"00001111",
"00001111",
"00111100",
"11110000",
"11000000",
"11000000",
"00000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00001111",
"00001111",
"11111111",
"11001111",
"11001111",
"11111100",
"00000000",
"00000000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11110000",
"11111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111100",
"00111100",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00001111",
"00001111",
"00001111",
"00001111",
"11111100",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00001111",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00001111",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00001111",
"00000011",
"00000000",
"00110000",
"11110000",
"00110000",
"00000000",
"00000000",
"00000011",
"00001111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00001111",
"00000011",
"00000000",
"00110000",
"11110000",
"00110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00001111",
"00001111",
"00000000",
"00000000",
"11111111",
"00001111",
"00001111",
"00001111",
"00111111",
"11110011",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"11111111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00001111",
"00111100",
"00111100",
"11110000",
"11110000",
"11110000",
"00111100",
"00111100",
"00001111",
"00001111",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00001111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00111111",
"11111111",
"11111111",
"11001111",
"11001111",
"11001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111100",
"11111100",
"11111100",
"11111100",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"11001111",
"11111111",
"11111100",
"11110000",
"00111100",
"00111111",
"00000000",
"00000000",
"11111100",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"11111100",
"11110000",
"00111100",
"00111100",
"00111100",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00001111",
"00001111",
"00000000",
"00000000",
"11111100",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11001111",
"11000011",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11110000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00001111",
"00001111",
"00001111",
"11001111",
"11001111",
"11001111",
"11001111",
"11001111",
"11111111",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"11110000",
"11110000",
"11000000",
"11000000",
"11000000",
"11000000",
"11110000",
"11110000",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00001111",
"00001111",
"00001111",
"00111111",
"11111100",
"11110000",
"11000000",
"11000000",
"11000000",
"11000000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00111100",
"11110000",
"11110000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00001100",
"00111100",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11110000",
"11110000",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11110000",
"00111100",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"11111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00111100",
"00111100",
"00111100",
"11111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00111100",
"11111100",
"00000000",
"00000000",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11001111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111100",
"00111100",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"00000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"00000000",
"11111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"11110000",
"11000000",
"11110000",
"00111100",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"11111111",
"11001111",
"11001111",
"11001111",
"00001111",
"00001111",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11001111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111100",
"00111100",
"00111100",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00001111",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00000000",
"00000000",
"11110000",
"00111100",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"00111100",
"00111100",
"11111100",
"11110000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00001111",
"11001111",
"11001111",
"11001111",
"11001111",
"11111111",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"11111100",
"11110000",
"11000000",
"11000000",
"11110000",
"11111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111100",
"11110000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00111100",
"11110000",
"11000000",
"00000000",
"00000000",
"00111100",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"11000000",
"11000000",
"11000000",
"11000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11111100",
"11111100",
"11000000",
"11000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11110000",
"00111100",
"00111100",
"00111100",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11110000",
"11111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111100",
"00111100",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00001111",
"00000011",
"00000000",
"00000000",
"11111100",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00001111",
"00001111",
"00001111",
"00001111",
"11111100",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00001111",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"11111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111111",
"00001111",
"00000000",
"00000000",
"00000000",
"11111111",
"00001111",
"00000011",
"00000000",
"00110000",
"11110000",
"00110000",
"00000000",
"00000000",
"00000011",
"00001111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"11000011",
"11000011",
"11000011",
"11000011",
"11001100",
"11110000",
"11001100",
"11000011",
"11000011",
"11000011",
"11000011",
"11000011",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00001111",
"00001111",
"00001111",
"00111100",
"11110000",
"00111100",
"00001111",
"00001111",
"00001111",
"00001111",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00001111",
"00111111",
"00111111",
"11111111",
"11001111",
"11001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00110000",
"11000000",
"00001111",
"00111111",
"00111111",
"11111111",
"11001111",
"11001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00001111",
"00111100",
"00111100",
"11110000",
"11110000",
"11110000",
"00111100",
"00111100",
"00001111",
"00001111",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00111111",
"11111111",
"11111111",
"11001111",
"11001111",
"11001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"11111111",
"00001111",
"00001111",
"00001111",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00001111",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"00001111",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11001111",
"11000011",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00111100",
"11110000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"00000000",
"11110000",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11110000",
"00000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"11110000",
"11110000",
"11000000",
"11000000",
"11000000",
"11000000",
"11110000",
"11110000",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111100",
"11111111",
"00001111",
"00000000",
"00000000",
"00000000",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"11111111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00001111",
"00001111",
"00001111",
"11001111",
"11001111",
"11001111",
"11001111",
"11001111",
"11001111",
"11001111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00001111",
"00001111",
"00001111",
"11001111",
"11001111",
"11001111",
"11001111",
"11001111",
"11001111",
"11001111",
"11111111",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00001111",
"00001111",
"00001111",
"00001111",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"11001111",
"11001111",
"11001111",
"11001111",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00001111",
"00001111",
"00001111",
"00001111",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00001111",
"00001111",
"00001111",
"00001111",
"11111111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"11001111",
"11001111",
"11001111",
"11001111",
"11001111",
"11001111",
"11001111",
"11001111",
"11001111",
"11001111",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"00000000",
"00000000",
"11110000",
"00111100",
"00111100",
"00111100",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11110000",
"11110000",
"11110000",
"00111100",
"00111100",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111100",
"00001100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00111100",
"00111100",
"11111100",
"00000000",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001100",
"00001100",
"00110000",
"11000000",
"11000000",
"00110000",
"00001100",
"00001100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00111100",
"11110000",
"00111100",
"00111100",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"00111100",
"00111100",
"11111100",
"11111100",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"00000000",
"00111100",
"00111100",
"00111100",
"00111100",
"11111100",
"11111100",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"11110000",
"11000000",
"11000000",
"11110000",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"11111100",
"11111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111100",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000011",
"00110000",
"00000011",
"00110000",
"00000011",
"00110000",
"00000011",
"00110000",
"00000011",
"00110000",
"00000011",
"00110000",
"00000011",
"00110000",
"00000011",
"00110000",
"00110011",
"11001100",
"00110011",
"11001100",
"00110011",
"11001100",
"00110011",
"11001100",
"00110011",
"11001100",
"00110011",
"11001100",
"00110011",
"11001100",
"00110011",
"11001100",
"11110011",
"00111111",
"11110011",
"00111111",
"11110011",
"00111111",
"11110011",
"00111111",
"11110011",
"00111111",
"11110011",
"00111111",
"11110011",
"00111111",
"11110011",
"00111111",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11111111",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"11000011",
"11000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"11111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11111111",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111111",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"00111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111111",
"11111111",
"00000000",
"00000000",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"00000000",
"00000000",
"11111111",
"11111111",
"11111111",
"11111111",
"00000000",
"00000000",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"00000000",
"00000000",
"11111111",
"11111111",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"00000011",
"00000011",
"11000011",
"11000011",
"11000011",
"11000011",
"11000011",
"11000011",
"11000011",
"11000011",
"00000011",
"00000011",
"11111111",
"11111111",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11000011",
"11000011",
"11000011",
"11000011",
"11000011",
"11000011",
"11000011",
"11000011",
"11000011",
"11000011",
"11000011",
"11000011",
"11000011",
"11000011",
"11000011",
"11000011",
"11110000",
"00111111",
"11110000",
"00000011",
"11110000",
"00111111",
"11110000",
"00000011",
"11110000",
"00111111",
"11110000",
"00000011",
"11110000",
"00111111",
"11110000",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"11111111",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"11111111",
"11111111",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00111100",
"00111100",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00111100",
"00000000",
"00000000",
"00111100",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"00111100",
"00111100",
"11110000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"00000000",
"11110000",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11110000",
"00000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"11110000",
"11000000",
"11000000",
"11110000",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111100",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"11111111",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00111100",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11110000",
"11110000",
"11110000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00111100",
"11111100",
"00111100",
"00111100",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00111100",
"00111100",
"00111100",
"11111100",
"00111100",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00000000",
"00000000",
"11111100",
"00000000",
"00000000",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11111100",
"11000000",
"11000000",
"00000000",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11110000",
"00111100",
"11110000",
"11000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11110000",
"00000000",
"00000000",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"11001111",
"11001111",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"00000000",
"11111100",
"00000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"11110000",
"00000000",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11110000",
"11110000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00000000",
"00000000",
"11000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"11000011",
"00110011",
"00000011",
"00000011",
"00110011",
"11000011",
"00001100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000"
	);

--------------------------------------------------------------------------
-- FONT hi byte
--------------------------------------------------------------------------
	signal RAM_FONT8_Hi: rom_type := (
--------------------------------------------------------------------------
-- FONT 8x8 1 bit on pixel
--------------------------------------------------------------------------
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",
"11110000",
"11110000",
"11110000",
"11110000",
"00001111",
"00001111",
"00001111",
"00001111",

--------------------------------------------------------------
---- FONT 8x8 2 bits on pixel
--------------------------------------------------------------
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00001100",
"00110011",
"00110000",
"00110011",
"00110000",
"00001100",
"00000011",
"00000011",
"00001111",
"00110000",
"00111111",
"00110000",
"00111100",
"00001111",
"00000011",
"00000000",
"00001111",
"00110000",
"00110000",
"00001100",
"00000011",
"00000000",
"00000000",
"00000000",
"00000011",
"00001100",
"00110000",
"00001100",
"00000011",
"00000000",
"00000000",
"00000000",
"00000011",
"00000000",
"00001100",
"00110011",
"00001100",
"00000000",
"00000011",
"00000000",
"00000011",
"00001100",
"00110000",
"00110000",
"00001111",
"00000000",
"00000011",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00111111",
"00111111",
"00111111",
"00111100",
"00111100",
"00111111",
"00111111",
"00111111",
"00000000",
"00000000",
"00000011",
"00001100",
"00001100",
"00000011",
"00000000",
"00000000",
"00111111",
"00111111",
"00111100",
"00110011",
"00110011",
"00111100",
"00111111",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00110000",
"00001111",
"00000000",
"00000011",
"00001100",
"00001100",
"00000011",
"00000000",
"00000000",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00001111",
"00000000",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00111111",
"00111111",
"00000000",
"00000000",
"00001100",
"00000011",
"00001111",
"00000011",
"00001100",
"00000000",
"00000000",
"00000000",
"00000000",
"00001100",
"00001111",
"00001111",
"00001111",
"00001100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00001111",
"00000011",
"00000011",
"00001111",
"00000011",
"00000000",
"00000000",
"00001100",
"00001100",
"00001100",
"00001100",
"00000000",
"00001100",
"00000000",
"00000000",
"00111111",
"11001100",
"00111100",
"00001100",
"00001100",
"00001100",
"00000000",
"00000000",
"00001111",
"00110000",
"00001111",
"00110000",
"00001111",
"00000000",
"00001111",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00001111",
"00000011",
"00000011",
"00001111",
"00000011",
"00111111",
"00000000",
"00000011",
"00001111",
"00000011",
"00000011",
"00000011",
"00000011",
"00000000",
"00000000",
"00000011",
"00000011",
"00000011",
"00000011",
"00001111",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00001100",
"00111111",
"00001100",
"00000011",
"00000000",
"00000000",
"00000000",
"00110000",
"00110000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110000",
"11111111",
"00110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00001111",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"00001111",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001100",
"00001100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001100",
"00111111",
"00001100",
"00111111",
"00001100",
"00000000",
"00000000",
"00000011",
"00111111",
"11000011",
"00111111",
"00000011",
"00111111",
"00000011",
"00000000",
"00111100",
"00111100",
"00000000",
"00000011",
"00001100",
"00110000",
"00000000",
"00000000",
"00000011",
"00001100",
"00000011",
"00001100",
"00110000",
"00001111",
"00000000",
"00000000",
"00000011",
"00000000",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000000",
"00000000",
"00110000",
"00001100",
"00111111",
"00001100",
"00110000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00111111",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000000",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00001100",
"00001100",
"00000000",
"00000000",
"00001111",
"00110000",
"00110000",
"00110011",
"00111100",
"00001111",
"00000000",
"00000000",
"00000000",
"00000011",
"00001100",
"00000000",
"00000000",
"00001111",
"00000000",
"00000000",
"00001111",
"00110000",
"00000000",
"00001111",
"00110000",
"00111111",
"00000000",
"00000000",
"00111111",
"00000000",
"00000000",
"00000000",
"00110000",
"00001111",
"00000000",
"00000000",
"00000000",
"00000011",
"00001100",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"00110000",
"00111111",
"00000000",
"00110000",
"00001111",
"00000000",
"00000000",
"00001111",
"00110000",
"00111111",
"00110000",
"00110000",
"00001111",
"00000000",
"00000000",
"00111111",
"00110000",
"00000000",
"00000000",
"00000011",
"00001100",
"00000000",
"00000000",
"00001111",
"00110000",
"00001111",
"00110000",
"00110000",
"00001111",
"00000000",
"00000000",
"00001111",
"00110000",
"00110000",
"00001111",
"00000000",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00000000",
"00000011",
"00000000",
"00000011",
"00000000",
"00000000",
"00000011",
"00001111",
"00111100",
"00001111",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"00000000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00000011",
"00000000",
"00000011",
"00001111",
"00000000",
"00000000",
"00001111",
"00110000",
"00000000",
"00000011",
"00000000",
"00000011",
"00000000",
"00001111",
"00110000",
"11000011",
"11001100",
"11001100",
"11000011",
"00110000",
"00001111",
"00000000",
"00000011",
"00001100",
"00110000",
"00111111",
"00110000",
"11111100",
"00000000",
"00000000",
"00111111",
"00001100",
"00001111",
"00001100",
"00001100",
"00111111",
"00000000",
"00000000",
"00001111",
"00110000",
"00110000",
"00110000",
"00110000",
"00001111",
"00000000",
"00000000",
"00111111",
"00001100",
"00001100",
"00001100",
"00001100",
"00111111",
"00000000",
"00000000",
"00111111",
"00001100",
"00001111",
"00001100",
"00001100",
"00111111",
"00000000",
"00000000",
"00111111",
"00001100",
"00001111",
"00001100",
"00001100",
"00111111",
"00000000",
"00000000",
"00001111",
"00110000",
"00110000",
"00110000",
"00110000",
"00001111",
"00000000",
"00000000",
"11111100",
"00110000",
"00111111",
"00110000",
"00110000",
"11111100",
"00000000",
"00000000",
"00111111",
"00000011",
"00000011",
"00000011",
"00000011",
"00111111",
"00000000",
"00000000",
"00001111",
"00000000",
"00000000",
"00000000",
"00110000",
"00001111",
"00000000",
"00000000",
"11111100",
"00110000",
"00111111",
"00110000",
"00110000",
"11111100",
"00000000",
"00000000",
"00110000",
"00110000",
"00110000",
"00110000",
"00110000",
"00111111",
"00000000",
"00000000",
"11110000",
"11110000",
"11001100",
"11000011",
"11000000",
"11110000",
"00000000",
"00000000",
"00110000",
"00111100",
"00110011",
"00110000",
"00110000",
"11110000",
"00000000",
"00000000",
"00001111",
"00110000",
"00110000",
"00110000",
"00110000",
"00001111",
"00000000",
"00000000",
"11111111",
"00110000",
"00110000",
"00111111",
"00110000",
"11111100",
"00000000",
"00000000",
"00001111",
"00110000",
"00110000",
"00110000",
"00110000",
"00001111",
"00000000",
"00000000",
"11111111",
"00110000",
"00110000",
"00111111",
"00110000",
"11111100",
"00000000",
"00000000",
"00001111",
"00110000",
"00001111",
"00000000",
"00110000",
"00001111",
"00000000",
"00000000",
"11111111",
"11000011",
"00000011",
"00000011",
"00000011",
"00001111",
"00000000",
"00000000",
"11111100",
"00110000",
"00110000",
"00110000",
"00110000",
"00001111",
"00000000",
"00000000",
"11110000",
"11000000",
"00110000",
"00110000",
"00001100",
"00000011",
"00000000",
"00000000",
"11110000",
"11000000",
"11000011",
"11000011",
"00111100",
"00110000",
"00000000",
"00000000",
"11110000",
"00001100",
"00000011",
"00001100",
"00110000",
"11110000",
"00000000",
"00000000",
"11110000",
"00110000",
"00001100",
"00000011",
"00000011",
"00001111",
"00000000",
"00000000",
"00111111",
"00110000",
"00000000",
"00000011",
"00001100",
"00111111",
"00000000",
"00000000",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000000",
"00000000",
"00001100",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00000000",
"00000000",
"00000000",
"00000011",
"00001100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00000000",
"00001111",
"00110000",
"00001111",
"00000000",
"00000000",
"00111100",
"00001100",
"00001111",
"00001100",
"00001100",
"00111111",
"00000000",
"00000000",
"00000000",
"00001111",
"00110000",
"00110000",
"00110000",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00110000",
"00110000",
"00001111",
"00000000",
"00000000",
"00000000",
"00001111",
"00110000",
"00111111",
"00110000",
"00001111",
"00000000",
"00000000",
"00000000",
"00000011",
"00001111",
"00000011",
"00000011",
"00001111",
"00000000",
"00000000",
"00000000",
"00001111",
"00110000",
"00110000",
"00001111",
"00000000",
"00001111",
"00000000",
"11110000",
"00110000",
"00111111",
"00110000",
"00110000",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000000",
"00000000",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000000",
"00000000",
"00110000",
"00001111",
"00000000",
"11110000",
"00110000",
"00110000",
"00111111",
"00110000",
"11111100",
"00000000",
"00000000",
"00001111",
"00000011",
"00000011",
"00000011",
"00000011",
"00001111",
"00000000",
"00000000",
"00000000",
"11001100",
"11110011",
"11000011",
"11000011",
"11000011",
"00000000",
"00000000",
"00000000",
"11110011",
"00111100",
"00110000",
"00110000",
"11111100",
"00000000",
"00000000",
"00000000",
"00001111",
"00110000",
"00110000",
"00110000",
"00001111",
"00000000",
"00000000",
"00000000",
"00111111",
"00001100",
"00001100",
"00001111",
"00001100",
"00111111",
"00000000",
"00000000",
"00001111",
"00110000",
"00110000",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00001111",
"00001100",
"00001100",
"00111111",
"00000000",
"00000000",
"00000000",
"00001111",
"00110000",
"00001111",
"00000000",
"00001111",
"00000000",
"00000000",
"00000011",
"00000011",
"00001111",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00110000",
"00110000",
"00110000",
"00001111",
"00000000",
"00000000",
"00000000",
"11111100",
"00110000",
"00001100",
"00001100",
"00000011",
"00000000",
"00000000",
"00000000",
"11110000",
"11000000",
"11000011",
"11001100",
"00110000",
"00000000",
"00000000",
"00000000",
"11111100",
"00001100",
"00000011",
"00001100",
"11111100",
"00000000",
"00000000",
"00000000",
"11110000",
"00001100",
"00001100",
"00000011",
"00000011",
"00111100",
"00000000",
"00000000",
"00111111",
"00000000",
"00000011",
"00001100",
"00111111",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00001111",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000000",
"00000000",
"00001111",
"00110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00001100",
"00111111",
"00000000",
"00000000",
"00001111",
"00110000",
"00110000",
"00111111",
"00110000",
"11110000",
"00000000",
"00000000",
"00111111",
"00001100",
"00001111",
"00001100",
"00001100",
"00111111",
"00000000",
"00000000",
"00111111",
"00001100",
"00001111",
"00001100",
"00001100",
"00111111",
"00000000",
"00000000",
"00001111",
"00000011",
"00000011",
"00000011",
"00000011",
"00001111",
"00000000",
"00000000",
"00000011",
"00001100",
"00001100",
"00001100",
"00001100",
"00111111",
"00110000",
"00000000",
"00111111",
"00001100",
"00001111",
"00001100",
"00001100",
"00111111",
"00000000",
"00000000",
"11110011",
"00110011",
"00001111",
"00110011",
"11000011",
"11000011",
"00000000",
"00000000",
"00001111",
"00110000",
"00000000",
"00000000",
"00110000",
"00001111",
"00000000",
"00000000",
"00110000",
"00110000",
"00110000",
"00110011",
"00111100",
"00110000",
"00000000",
"00000011",
"00110000",
"00110000",
"00110000",
"00110011",
"00111100",
"00110000",
"00000000",
"00000000",
"00111100",
"00001100",
"00001111",
"00001100",
"00001100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000011",
"00001100",
"00001100",
"00001100",
"00111100",
"00000000",
"00000000",
"11110000",
"00111100",
"00110011",
"00110011",
"00110000",
"11111100",
"00000000",
"00000000",
"11111100",
"00110000",
"00111111",
"00110000",
"00110000",
"11111100",
"00000000",
"00000000",
"00001111",
"00110000",
"00110000",
"00110000",
"00110000",
"00001111",
"00000000",
"00000000",
"11111111",
"00110000",
"00110000",
"00110000",
"00110000",
"11111100",
"00000000",
"00000000",
"00111111",
"00001100",
"00001100",
"00001111",
"00001100",
"00111111",
"00000000",
"00000000",
"00001111",
"00110000",
"00110000",
"00110000",
"00110000",
"00001111",
"00000000",
"00000000",
"00111111",
"00110011",
"00000011",
"00000011",
"00000011",
"00001111",
"00000000",
"00000000",
"11110000",
"00110000",
"00001100",
"00000011",
"00000000",
"00111111",
"00000000",
"00000000",
"00000011",
"00111111",
"11000011",
"11000011",
"11000011",
"00111111",
"00000011",
"00000000",
"00111100",
"00001100",
"00000011",
"00000011",
"00001100",
"00111100",
"00000000",
"00000000",
"11111100",
"00110000",
"00110000",
"00110000",
"00110000",
"11111111",
"00000000",
"00000000",
"11111100",
"00110000",
"00110000",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"11000011",
"11000011",
"11000011",
"11000011",
"11000011",
"11111111",
"00000000",
"00000000",
"11000011",
"11000011",
"11000011",
"11000011",
"11000011",
"11111111",
"00000000",
"00000000",
"11111100",
"11001100",
"00001111",
"00001100",
"00001100",
"00111111",
"00000000",
"00000000",
"11111100",
"00110000",
"00111111",
"00110000",
"00110000",
"11111111",
"00000000",
"00000000",
"00111111",
"00001100",
"00001111",
"00001100",
"00001100",
"00111111",
"00000000",
"00000000",
"00001111",
"00110000",
"00000011",
"00000000",
"00110000",
"00001111",
"00000000",
"00000000",
"11000011",
"11001100",
"11001100",
"11111100",
"11001100",
"11000011",
"00000000",
"00000000",
"00001111",
"00110000",
"00110000",
"00001111",
"00000011",
"00111100",
"00000000",
"00000000",
"00000000",
"00001111",
"00000000",
"00001111",
"00110000",
"00001111",
"00000000",
"00000000",
"00001111",
"00110000",
"00001111",
"00110000",
"00110000",
"00001111",
"00000000",
"00000000",
"00000000",
"00111111",
"00001100",
"00001111",
"00001100",
"00111111",
"00000000",
"00000000",
"00000000",
"00111111",
"00001100",
"00001100",
"00001100",
"00111111",
"00000000",
"00000000",
"00000000",
"00001111",
"00000011",
"00001100",
"00001100",
"00111111",
"00110000",
"00000000",
"00000000",
"00001111",
"00110000",
"00111111",
"00110000",
"00001111",
"00000000",
"00000000",
"00000000",
"11110011",
"00110011",
"00001111",
"00110011",
"11110011",
"00000000",
"00000000",
"00000000",
"00001111",
"00110000",
"00000000",
"00110000",
"00001111",
"00000000",
"00000000",
"00000000",
"11111100",
"00110000",
"00110000",
"00110011",
"11111100",
"00000000",
"00000011",
"00000000",
"11111100",
"00110000",
"00110000",
"00110011",
"11111100",
"00000000",
"00000000",
"00000000",
"11111100",
"00110000",
"00111111",
"00110000",
"11111100",
"00000000",
"00000000",
"00000000",
"00001111",
"00000011",
"00000011",
"00001100",
"00111100",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11001100",
"11000011",
"11000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00110000",
"00111111",
"00110000",
"11111100",
"00000000",
"00000000",
"00000000",
"00001111",
"00110000",
"00110000",
"00110000",
"00001111",
"00000000",
"00000000",
"00000000",
"11111111",
"00110000",
"00110000",
"00110000",
"11111100",
"00000000",
"11000000",
"00001100",
"11000000",
"00001100",
"11000000",
"00001100",
"11000000",
"00001100",
"11000011",
"00110000",
"11000011",
"00110000",
"11000011",
"00110000",
"11000011",
"00000000",
"11001100",
"00110011",
"11001100",
"00110011",
"11001100",
"00110011",
"11001100",
"00000000",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"11111111",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"11111111",
"00000011",
"11111111",
"00000011",
"00000011",
"00000011",
"00001100",
"00001100",
"00001100",
"11111100",
"00001100",
"00001100",
"00001100",
"00001100",
"00000000",
"00000000",
"00000000",
"11111111",
"00001100",
"00001100",
"00001100",
"00001100",
"00000000",
"00000000",
"11111111",
"00000011",
"11111111",
"00000011",
"00000011",
"00000011",
"00001100",
"00001100",
"11111100",
"00000000",
"11111100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00000000",
"00000000",
"11111111",
"00000000",
"11111100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"11111100",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00001100",
"00001100",
"00001100",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"11111111",
"00000011",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00000011",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00000011",
"11111111",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"11111100",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"11111100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00000000",
"00000000",
"11111111",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00001100",
"00001100",
"11111100",
"00000000",
"11111100",
"00001100",
"00001100",
"00001100",
"00000011",
"00000011",
"11111111",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00001100",
"00001100",
"00001100",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"11111111",
"00000011",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"11111111",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00001111",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"00001100",
"11111100",
"00001100",
"00001100",
"00001100",
"00001100",
"00000011",
"00000011",
"11111111",
"00000000",
"11111111",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"00001100",
"00001100",
"00001111",
"00001100",
"00111111",
"00000000",
"00000000",
"00001111",
"00110000",
"00110000",
"00110000",
"00001111",
"00000000",
"00000000",
"00000000",
"00111111",
"00110011",
"00000011",
"00000011",
"00001111",
"00000000",
"00000000",
"00000000",
"11111100",
"00110000",
"00110000",
"00001111",
"00000000",
"00111111",
"00000000",
"00000000",
"00000011",
"00111111",
"11000011",
"11000011",
"00111111",
"00000011",
"00000000",
"00000000",
"11111100",
"00001100",
"00000011",
"00001100",
"11111100",
"00000000",
"00000000",
"00000000",
"11111100",
"00110000",
"00110000",
"00110000",
"11111111",
"00000000",
"00000000",
"00000000",
"11111100",
"00110000",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000011",
"11000011",
"11000011",
"11000011",
"11111111",
"00000000",
"00000000",
"00000000",
"11000011",
"11000011",
"11000011",
"11000011",
"11111111",
"00000000",
"00000000",
"00000000",
"11111100",
"11001100",
"00001111",
"00001100",
"00111111",
"00000000",
"00000000",
"00000000",
"11111100",
"00110000",
"00111111",
"00110000",
"11111111",
"00000000",
"00000000",
"00000000",
"00111111",
"00001100",
"00001111",
"00001100",
"00111111",
"00000000",
"00000000",
"00000000",
"00001111",
"00110000",
"00000011",
"00110000",
"00001111",
"00000000",
"00000000",
"00000000",
"11000011",
"11001100",
"11111100",
"11001100",
"11000011",
"00000000",
"00000000",
"00000000",
"00001111",
"00110000",
"00001111",
"00001100",
"00111100",
"00000000",
"00001100",
"00111111",
"00001100",
"00001111",
"00001100",
"00001100",
"00111111",
"00000000",
"00001100",
"00000000",
"00001111",
"00110000",
"00111111",
"00110000",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00001111",
"00000011",
"00000011",
"00001111",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00001100",
"00111111",
"00001100",
"00000011",
"00000000",
"00000000",
"00000011",
"00001111",
"00110011",
"00000011",
"00000011",
"00000011",
"00000000",
"00000000",
"00000011",
"00000011",
"00000011",
"00110011",
"00001111",
"00000011",
"00000000",
"00000000",
"00000011",
"00000000",
"00111111",
"00000000",
"00000011",
"00000000",
"00000000",
"00000011",
"00000011",
"00111111",
"00000011",
"00000011",
"00000000",
"00111111",
"00000000",
"00000000",
"11000000",
"11000000",
"11110000",
"11001100",
"11000011",
"11000000",
"00000000",
"00000000",
"00000000",
"00110000",
"00001111",
"00110000",
"00001111",
"00110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000"
);

--------------------------------------------------------------
--
--------------------------------------------------------------

	signal RAM_FONT16_Hi: rom_type := (
--------------------------------------------------------------
---- FONT 16x16 1 bit on pixel or 8x16 2 bits on pixel
--------------------------------------------------------------
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"11000000",
"11001100",
"11000000",
"11000000",
"11001111",
"11000011",
"11000000",
"11000000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"11111111",
"11110011",
"11111111",
"11111111",
"11110000",
"11111100",
"11111111",
"11111111",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110000",
"11110000",
"00110000",
"00110000",
"00110000",
"00000011",
"00001100",
"00110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110000",
"11110000",
"00110000",
"00110000",
"00110000",
"00000011",
"00001100",
"00110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00001111",
"00001111",
"00000011",
"00111100",
"11111111",
"11111111",
"00111100",
"00000011",
"00001111",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00001111",
"00001111",
"00111111",
"11111111",
"11111111",
"11111111",
"00111111",
"00000011",
"00001111",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00001111",
"00001111",
"00001111",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"11111111",
"11111111",
"11111100",
"11110000",
"11110000",
"11110000",
"11111100",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00001111",
"00111100",
"00110000",
"00110000",
"00110000",
"00111100",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"11111111",
"11110000",
"11000011",
"11001111",
"11001111",
"11001111",
"11000011",
"11110000",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"00000000",
"00000011",
"00000000",
"00000011",
"00001111",
"00111111",
"11110000",
"11110000",
"11110000",
"11110000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00111100",
"00111100",
"00111100",
"00111100",
"00001111",
"00000011",
"00111111",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00111111",
"11111111",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"00111100",
"00111100",
"00111111",
"00111100",
"00111100",
"00111100",
"00111100",
"11111100",
"11111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"11110011",
"00001111",
"11111100",
"11111100",
"00001111",
"11110011",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11110000",
"11111100",
"11111111",
"11111111",
"11111111",
"11111111",
"11111100",
"11110000",
"11000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"11111111",
"11111111",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00001111",
"00111111",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00111111",
"00001111",
"00000011",
"00000000",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00000000",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"11110011",
"11110011",
"11110011",
"11110011",
"11110011",
"00111111",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"11110000",
"00111100",
"00001111",
"00111100",
"11110000",
"11110000",
"00111100",
"00001111",
"00000000",
"11110000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00001111",
"00111111",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00111111",
"00001111",
"00000011",
"00111111",
"00000000",
"00000000",
"00000000",
"00000011",
"00001111",
"00111111",
"11111111",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"11111111",
"00111111",
"00001111",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00001111",
"00111111",
"11111111",
"00111111",
"00001111",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001100",
"00111100",
"11111111",
"00111100",
"00001100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00001111",
"00001111",
"00111111",
"00111111",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"00111111",
"00111111",
"00001111",
"00001111",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00001111",
"00111111",
"00111111",
"00111111",
"00111111",
"00001111",
"00000011",
"00000011",
"00000000",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"00111100",
"11111111",
"11111111",
"00111100",
"00111100",
"00111100",
"11111111",
"11111111",
"00111100",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00111111",
"11110011",
"11110011",
"11110011",
"11110011",
"00111111",
"00000011",
"00000011",
"11110011",
"11110011",
"00111111",
"00000011",
"00000011",
"00000000",
"00000000",
"11111100",
"11001100",
"11111100",
"00000000",
"00000011",
"00000011",
"00001111",
"00001111",
"00111100",
"00111100",
"11110000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00111100",
"00111100",
"00111100",
"00001111",
"00111111",
"11110011",
"11110011",
"11110000",
"11110000",
"11110000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00001111",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"00001111",
"11111111",
"11111111",
"00001111",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00111111",
"00111111",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00001111",
"00001111",
"00111100",
"00111100",
"11110000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"11110000",
"11110000",
"11110000",
"11110000",
"11110011",
"11110011",
"11111100",
"11111100",
"11110000",
"11110000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000010",
"00001010",
"00101010",
"00000010",
"00000010",
"00000010",
"00000010",
"00000010",
"00000010",
"00000010",
"00000010",
"00101010",
"00000000",
"00000000",
"00000000",
"00000000",
"00000101",
"00010100",
"01010000",
"01010000",
"00000000",
"00000000",
"00000000",
"00000001",
"00000101",
"00010100",
"01010000",
"01010101",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11110000",
"00000000",
"00000011",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00001111",
"00001111",
"00111100",
"00111100",
"11110000",
"11110000",
"11111111",
"00000000",
"00000000",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11110000",
"11110000",
"11110000",
"11111111",
"11111100",
"11110000",
"00000000",
"00000000",
"11110000",
"00111100",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00111100",
"11110000",
"11110000",
"11111111",
"11111100",
"11110000",
"11110000",
"11110000",
"11110000",
"00111100",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11110000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00111100",
"11110000",
"11110000",
"00111100",
"00001111",
"00111100",
"11110000",
"11110000",
"11110000",
"00111100",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00111100",
"11110000",
"11110000",
"11110000",
"11110000",
"00111100",
"00001111",
"00000000",
"00111100",
"00111100",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00001111",
"00111111",
"00001111",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"00111111",
"00000000",
"00111111",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"00111100",
"00001111",
"00000011",
"00000000",
"00000000",
"00000000",
"00000011",
"00001111",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00111100",
"11110000",
"11110000",
"11110000",
"00000000",
"00000000",
"00000011",
"00000011",
"00000000",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"11110000",
"11110000",
"11110011",
"11110011",
"11110011",
"11110011",
"11110000",
"11110000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00001111",
"00111111",
"11111100",
"11110000",
"11110000",
"11110000",
"11110000",
"11111111",
"11110000",
"11110000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00111100",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00111100",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00111100",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00111100",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11111111",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11111100",
"11111111",
"11111111",
"11110011",
"11110011",
"11110011",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11111100",
"11111100",
"11111111",
"11111111",
"11110011",
"11110011",
"11110000",
"11110000",
"11110000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00111100",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00111100",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111111",
"00111100",
"00111100",
"00111100",
"00111100",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00111100",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00111111",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111111",
"00111100",
"00111100",
"00111100",
"00111100",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"11110000",
"11110000",
"11110000",
"11110000",
"00111111",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11110011",
"11000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00111111",
"00001111",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110011",
"11110011",
"11110011",
"11110011",
"11110011",
"11111111",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"00111100",
"00111100",
"00001111",
"00001111",
"00001111",
"00001111",
"00111100",
"00111100",
"11110000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11111100",
"00111111",
"00001111",
"00000011",
"00000011",
"00000011",
"00000011",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11110000",
"11000000",
"00000000",
"00000011",
"00000011",
"00001111",
"00001111",
"00111100",
"00111100",
"11110000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"00111100",
"00111100",
"00001111",
"00001111",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00001111",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"00000000",
"00000000",
"00001111",
"00001111",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00000000",
"00001111",
"00111100",
"00111100",
"00111100",
"00111100",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00111100",
"00111100",
"00111100",
"00111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11110011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"11110000",
"11110000",
"11111111",
"11110000",
"11110000",
"11110000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00111100",
"00111100",
"00111100",
"11111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00111111",
"00000000",
"11110000",
"00111111",
"00000000",
"11111100",
"00111100",
"00111100",
"00111100",
"00111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00000000",
"00001111",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00111100",
"00001111",
"00000000",
"11111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111111",
"00111100",
"00111100",
"00111100",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"11111111",
"11110011",
"11110011",
"11110011",
"11110000",
"11110000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110011",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110011",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111111",
"00111100",
"00111100",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110011",
"00111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"11110000",
"11110000",
"00111111",
"00000011",
"00000000",
"11110000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00001111",
"00001111",
"11111111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11111100",
"00111111",
"00001111",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110011",
"11110011",
"11110011",
"11110011",
"11111111",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11111100",
"00111111",
"00001111",
"00001111",
"00111111",
"11111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00111111",
"00000000",
"00000011",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11110000",
"00000000",
"00000011",
"00001111",
"00111100",
"11110000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00000011",
"00000011",
"00111111",
"00111111",
"00000011",
"00000011",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000000",
"00000000",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"11110011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00001111",
"00111100",
"11110000",
"11110000",
"11110000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00001111",
"00111111",
"11111100",
"11110000",
"11110000",
"11110000",
"11110000",
"11111111",
"11110000",
"11110000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00001111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111111",
"11110000",
"00000000",
"00000000",
"00000000",
"11111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"11000011",
"11000011",
"11000011",
"11000011",
"00110011",
"00001111",
"00110011",
"11000011",
"11000011",
"11000011",
"11000011",
"11000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"11110000",
"11110000",
"00000000",
"00000000",
"00000011",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110011",
"11110011",
"11111111",
"11111100",
"11111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001100",
"00000011",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110011",
"11110011",
"11111111",
"11111100",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11111100",
"11111111",
"11111111",
"11110011",
"11110011",
"11110011",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11111111",
"11110000",
"11110000",
"11110000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00111100",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00111100",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111111",
"00111100",
"00111100",
"00111100",
"00111100",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00111100",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00111100",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11110011",
"11000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00111100",
"00001111",
"00000011",
"00111111",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00000011",
"00111111",
"11110011",
"11110011",
"11110011",
"11110011",
"11110011",
"11110011",
"00111111",
"00000011",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"00111100",
"00111100",
"00001111",
"00001111",
"00001111",
"00001111",
"00111100",
"00111100",
"11110000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110011",
"11110011",
"11110011",
"11110011",
"11110011",
"11110011",
"11110011",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110011",
"11110011",
"11110011",
"11110011",
"11110011",
"11110011",
"11110011",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11111111",
"11110011",
"11110011",
"11110011",
"11110011",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11111111",
"11110000",
"11110000",
"11110000",
"11110000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"11110000",
"11110000",
"00000000",
"00000000",
"00000011",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110011",
"11110011",
"11110011",
"11110011",
"11111111",
"11111111",
"11110011",
"11110011",
"11110011",
"11110011",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00111111",
"00001111",
"00111100",
"00111100",
"00111100",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"11110000",
"00000000",
"00111111",
"11110000",
"11110000",
"11110000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00111100",
"11110000",
"11111111",
"11110000",
"11110000",
"11110000",
"11110000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11110000",
"11110000",
"11111111",
"11110000",
"11110000",
"11110000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00111100",
"00111100",
"00111100",
"00111100",
"11110000",
"11111111",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"11110000",
"11110000",
"11110000",
"11111111",
"11110000",
"11110000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000011",
"11000011",
"00110011",
"00001111",
"00001111",
"00110011",
"11000011",
"11000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"11110000",
"11110000",
"00000011",
"00000000",
"11110000",
"11110000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110011",
"11111111",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001100",
"00000011",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110011",
"11111111",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11111111",
"11111111",
"11110000",
"11110000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11111100",
"11111111",
"11110011",
"11110011",
"11110000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11111111",
"11110000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000011",
"00110000",
"00000011",
"00110000",
"00000011",
"00110000",
"00000011",
"00110000",
"00000011",
"00110000",
"00000011",
"00110000",
"00000011",
"00110000",
"00000011",
"00110000",
"00110011",
"11001100",
"00110011",
"11001100",
"00110011",
"11001100",
"00110011",
"11001100",
"00110011",
"11001100",
"00110011",
"11001100",
"00110011",
"11001100",
"00110011",
"11001100",
"11110011",
"00111111",
"11110011",
"00111111",
"11110011",
"00111111",
"11110011",
"00111111",
"11110011",
"00111111",
"11110011",
"00111111",
"11110011",
"00111111",
"11110011",
"00111111",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"11111111",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"11111111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000011",
"11111111",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"11111111",
"00000000",
"11111111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"11111111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"11111111",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"11111111",
"00000011",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000011",
"11000011",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11000000",
"11111111",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"11111111",
"11111111",
"00000000",
"00000000",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"00000000",
"00000000",
"11111111",
"11111111",
"11111111",
"11111111",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11111111",
"11111111",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"00000000",
"00000000",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"00000000",
"00000000",
"11111111",
"11111111",
"11111111",
"11111111",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11111111",
"11111111",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"00001111",
"11000000",
"00001111",
"11111100",
"00001111",
"11000000",
"00001111",
"11111100",
"00001111",
"11000000",
"00001111",
"11111100",
"00001111",
"11000000",
"00001111",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11111111",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11111111",
"11111111",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11111111",
"11111111",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11110000",
"11110000",
"11110000",
"11110000",
"11111111",
"11110000",
"11110000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11110000",
"00111100",
"00001111",
"00001111",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00000011",
"00111111",
"11110011",
"11110011",
"11110011",
"11110011",
"11110011",
"00111111",
"00000011",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"00111100",
"00001111",
"00001111",
"00111100",
"11110000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11110000",
"11110000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11000011",
"11000011",
"11000011",
"11000011",
"11000011",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000000",
"11000000",
"11000011",
"11000011",
"11000011",
"11000011",
"11000011",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11001111",
"11001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11111100",
"11110011",
"11110011",
"11110011",
"11111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11110000",
"11110000",
"11110000",
"11111111",
"11110000",
"11110000",
"11110000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"11000000",
"11000000",
"00000011",
"00000000",
"11000000",
"11000000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11000011",
"11001111",
"11001111",
"11001111",
"11111111",
"11001111",
"11001111",
"11000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"11110000",
"11110000",
"11110000",
"00111111",
"00001111",
"00111100",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"00000000",
"11111111",
"00000000",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00111111",
"00000011",
"00000011",
"00000000",
"00000000",
"11111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00000011",
"00000000",
"00000000",
"00000000",
"00000011",
"00001111",
"00000000",
"00000000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00001111",
"00111100",
"00001111",
"00000011",
"00000000",
"00000000",
"00000000",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"00000011",
"11110011",
"11110011",
"11110011",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00000000",
"00111111",
"00000000",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"11110011",
"00000000",
"00111111",
"11110011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00111100",
"00111100",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111100",
"00111100",
"00111100",
"00111100",
"00001111",
"00000011",
"00000000",
"00000000",
"11110011",
"00111100",
"00111100",
"00111100",
"00111100",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001111",
"00110000",
"11000011",
"11001100",
"11001100",
"11001100",
"11001100",
"11000011",
"00110000",
"00001111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111111",
"00111111",
"00111111",
"00111111",
"00111111",
"00111111",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000"
	);

--------------------------------------------------------------------------
-- COLOR Table
--------------------------------------------------------------------------
	type rem_type is array (0 to 255) of std_logic_vector(7 downto 0);
	signal RAM_COLOR_Lo: rem_type := (
x"03",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",
x"03",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",
x"03",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",
x"03",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",
x"03",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",
x"03",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",
x"03",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",
x"03",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",
x"03",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",
x"03",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",
x"03",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",
x"03",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",
x"03",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",
x"03",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",
x"03",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",
x"03",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF"
	);

	signal RAM_COLOR_Hi: rem_type := (
x"7F",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",
x"7F",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",
x"7F",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",
x"7F",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",
x"7F",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",
x"7F",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",
x"7F",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",
x"7F",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",
x"7F",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",
x"7F",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",
x"7F",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",
x"7F",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",
x"7F",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",
x"7F",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",
x"7F",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",
x"7F",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01",x"23",x"45",x"67",x"89",x"AB",x"CD",x"EF",x"01"
	);

begin

process (clk)
begin
  if rising_edge(clk) then

    if ( addr_r(15) = '0' ) then
        data_r( 7 downto 0) <= RAM_SCREEN_Lo(to_integer(unsigned(addr_r(14 downto 0))));
        data_r(15 downto 8) <= RAM_SCREEN_Hi(to_integer(unsigned(addr_r(14 downto 0))));
    else
      if ( addr_r(15 downto 8) = "11111111" ) then
          data_r( 7 downto 0) <= RAM_COLOR_Lo(to_integer(unsigned(addr_r(7 downto 0))));
          data_r(15 downto 8) <= RAM_COLOR_Hi(to_integer(unsigned(addr_r(7 downto 0))));
      else
        if ( addr_r(14 downto 13) = "11" ) then
          data_r( 7 downto 0) <= RAM_FONT8_Lo(to_integer(unsigned(addr_r(12 downto 0))));
          data_r(15 downto 8) <= RAM_FONT8_Hi(to_integer(unsigned(addr_r(12 downto 0))));
        else
          data_r( 7 downto 0) <= RAM_FONT16_Lo(to_integer(unsigned(addr_r(12 downto 0))));
          data_r(15 downto 8) <= RAM_FONT16_Hi(to_integer(unsigned(addr_r(12 downto 0))));
--        elsif ( addr_r(14 downto 13) = "11" ) then
        end if;
      end if;
    end if;

    if ( we = '0' ) then
      if ( addr_w(15) = '0' ) then
        if ( le = '0' ) then
          RAM_SCREEN_Lo(to_integer(unsigned(addr_w(14 downto 0)))) <= data_w( 7 downto 0);
        end if;
        if ( he = '0' ) then
          RAM_SCREEN_Hi(to_integer(unsigned(addr_w(14 downto 0)))) <= data_w(15 downto 8);
        end if;
      else
        if ( addr_r(15 downto 8) = "11111111" ) then
          if ( le = '0' ) then
            RAM_COLOR_Lo(to_integer(unsigned(addr_w(7 downto 0)))) <= data_w( 7 downto 0);
          end if;
          if ( he = '0' ) then
            RAM_COLOR_Hi(to_integer(unsigned(addr_w(7 downto 0)))) <= data_w(15 downto 8);
          end if;
        else
          if ( addr_r(14 downto 13) = "11" ) then
            if ( le = '0' ) then
              RAM_FONT8_Lo(to_integer(unsigned(addr_w(12 downto 0)))) <= data_w( 7 downto 0);
            end if;
            if ( he = '0' ) then
              RAM_FONT8_Hi(to_integer(unsigned(addr_w(12 downto 0)))) <= data_w(15 downto 8);
            end if;
          else
            if ( le = '0' ) then
              RAM_FONT16_Lo(to_integer(unsigned(addr_w(12 downto 0)))) <= data_w( 7 downto 0);
            end if;
            if ( he = '0' ) then
              RAM_FONT16_Hi(to_integer(unsigned(addr_w(12 downto 0)))) <= data_w(15 downto 8);
            end if;
          end if;
        end if;
      end if;
    end if;

  end if;

end process;
	
end Behavioral;