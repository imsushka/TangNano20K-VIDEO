LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY mapper IS 
	PORT
	(
		RESET_n :  IN  STD_LOGIC;
		CLK   :  IN  STD_LOGIC;

		A     :  IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		D     :  IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		WR    :  IN  STD_LOGIC;

		Q     :  OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
		SET   :  OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END mapper;

ARCHITECTURE bdf_type OF mapper IS 

SIGNAL	Q_ALT :   STD_LOGIC_VECTOR(11 DOWNTO 0);
SIGNAL	SET_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SET_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SET_2 : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SET_3 : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SET_4 : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SET_5 : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SET_6 : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SET_7 : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	W :       STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	DFF_0 :   STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	DFF_1 :   STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	DFF_2 :   STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	DFF_3 :   STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	DFF_4 :   STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	DFF_5 :   STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	DFF_6 :   STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	DFF_7 :   STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	DFF_8 :   STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	DFF_9 :   STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	DFF_A :   STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	DFF_B :   STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	DFF_C :   STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	DFF_D :   STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	DFF_E :   STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	DFF_F :   STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	ABUF :    STD_LOGIC_VECTOR(2 DOWNTO 0);

SIGNAL	EQ :      STD_LOGIC;
SIGNAL	EQ0 :     STD_LOGIC;
SIGNAL	EQ1 :     STD_LOGIC;
SIGNAL	EQ2 :     STD_LOGIC;
SIGNAL	EQ3 :     STD_LOGIC;
SIGNAL	EQ4 :     STD_LOGIC;
SIGNAL	EQ5 :     STD_LOGIC;
SIGNAL	EQ6 :     STD_LOGIC;
SIGNAL	EQ7 :     STD_LOGIC;
SIGNAL	WR00 :    STD_LOGIC;
SIGNAL	WR01 :    STD_LOGIC;
SIGNAL	WR10 :    STD_LOGIC;
SIGNAL	WR11 :    STD_LOGIC;
SIGNAL	WR20 :    STD_LOGIC;
SIGNAL	WR21 :    STD_LOGIC;
SIGNAL	WR30 :    STD_LOGIC;
SIGNAL	WR31 :    STD_LOGIC;
SIGNAL	WR40 :    STD_LOGIC;
SIGNAL	WR41 :    STD_LOGIC;
SIGNAL	WR50 :    STD_LOGIC;
SIGNAL	WR51 :    STD_LOGIC;
SIGNAL	WR60 :    STD_LOGIC;
SIGNAL	WR61 :    STD_LOGIC;
SIGNAL	WR70 :    STD_LOGIC;
SIGNAL	WR71 :    STD_LOGIC;

BEGIN 

EQ  <= '1' WHEN A(2 DOWNTO 0) = ABUF  ELSE '0';

EQ0 <= '1' WHEN A(2 DOWNTO 0) = "000" ELSE '0';
EQ1 <= '1' WHEN A(2 DOWNTO 0) = "001" ELSE '0';
EQ2 <= '1' WHEN A(2 DOWNTO 0) = "010" ELSE '0';
EQ3 <= '1' WHEN A(2 DOWNTO 0) = "011" ELSE '0';
EQ4 <= '1' WHEN A(2 DOWNTO 0) = "100" ELSE '0';
EQ5 <= '1' WHEN A(2 DOWNTO 0) = "101" ELSE '0';
EQ6 <= '1' WHEN A(2 DOWNTO 0) = "110" ELSE '0';
EQ7 <= '1' WHEN A(2 DOWNTO 0) = "111" ELSE '0';

WR00 <= NOT(EQ) AND EQ0 AND NOT(WR);
WR01 <=     EQ  AND EQ0 AND NOT(WR);
WR10 <= NOT(EQ) AND EQ1 AND NOT(WR);
WR11 <=     EQ  AND EQ1 AND NOT(WR);
WR20 <= NOT(EQ) AND EQ2 AND NOT(WR);
WR21 <=     EQ  AND EQ2 AND NOT(WR);
WR30 <= NOT(EQ) AND EQ3 AND NOT(WR);
WR31 <=     EQ  AND EQ3 AND NOT(WR);
WR40 <= NOT(EQ) AND EQ4 AND NOT(WR);
WR41 <=     EQ  AND EQ4 AND NOT(WR);
WR50 <= NOT(EQ) AND EQ5 AND NOT(WR);
WR51 <=     EQ  AND EQ5 AND NOT(WR);
WR60 <= NOT(EQ) AND EQ6 AND NOT(WR);
WR61 <=     EQ  AND EQ6 AND NOT(WR);
WR70 <= NOT(EQ) AND EQ7 AND NOT(WR);
WR71 <=     EQ  AND EQ7 AND NOT(WR);

PROCESS(WR)
BEGIN
  IF ( RISING_EDGE(WR) ) THEN
    ABUF <= A(2 DOWNTO 0);
  END IF;
END PROCESS;

PROCESS(WR00, RESET_n)
BEGIN
  IF (RESET_n = '0') THEN
    DFF_0 <= "11111111";
  ELSIF (FALLING_EDGE(WR00)) THEN
    DFF_0 <= D;
  END IF;
END PROCESS;

PROCESS(WR01, RESET_n)
BEGIN
  IF (RESET_n = '0') THEN
    DFF_8 <= "1111";
    SET_0 <= "1111";
  ELSIF (FALLING_EDGE(WR01)) THEN
    DFF_8 <= D(3 DOWNTO 0);
    SET_0 <= D(7 DOWNTO 4);
  END IF;
END PROCESS;

PROCESS(WR10, RESET_n)
BEGIN
  IF (RESET_n = '0') THEN
    DFF_1 <= "11111111";
  ELSIF (FALLING_EDGE(WR10)) THEN
    DFF_1 <= D;
  END IF;
END PROCESS;

PROCESS(WR11, RESET_n)
BEGIN
  IF (RESET_n = '0') THEN
    DFF_9 <= "1111";
    SET_1 <= "1111";
  ELSIF (FALLING_EDGE(WR11)) THEN
    DFF_9 <= D(3 DOWNTO 0);
    SET_1 <= D(7 DOWNTO 4);
  END IF;
END PROCESS;

PROCESS(WR20, RESET_n)
BEGIN
  IF (RESET_n = '0') THEN
    DFF_2 <= "11111111";
  ELSIF (FALLING_EDGE(WR20)) THEN
    DFF_2 <= D;
  END IF;
END PROCESS;

PROCESS(WR21, RESET_n)
BEGIN
  IF (RESET_n = '0') THEN
    DFF_A <= "1111";
    SET_2 <= "1111";
  ELSIF (FALLING_EDGE(WR21)) THEN
    DFF_A <= D(3 DOWNTO 0);
    SET_2 <= D(7 DOWNTO 4);
  END IF;
END PROCESS;

PROCESS(WR30, RESET_n)
BEGIN
  IF (RESET_n = '0') THEN
    DFF_3 <= "11111111";
  ELSIF (FALLING_EDGE(WR30)) THEN
    DFF_3 <= D;
  END IF;
END PROCESS;

PROCESS(WR31, RESET_n)
BEGIN
  IF (RESET_n = '0') THEN
    DFF_B <= "1111";
    SET_3 <= "1111";
  ELSIF (FALLING_EDGE(WR31)) THEN
    DFF_B <= D(3 DOWNTO 0);
    SET_3 <= D(7 DOWNTO 4);
  END IF;
END PROCESS;

PROCESS(WR40, RESET_n)
BEGIN
  IF (RESET_n = '0') THEN
    DFF_4 <= "11111111";
  ELSIF (FALLING_EDGE(WR40)) THEN
    DFF_4 <= D;
  END IF;
END PROCESS;

PROCESS(WR41, RESET_n)
BEGIN
  IF (RESET_n = '0') THEN
    DFF_C <= "1111";
    SET_4 <= "1111";
  ELSIF (FALLING_EDGE(WR41)) THEN
    DFF_C <= D(3 DOWNTO 0);
    SET_4 <= D(7 DOWNTO 4);
  END IF;
END PROCESS;

PROCESS(WR50, RESET_n)
BEGIN
  IF (RESET_n = '0') THEN
    DFF_5 <= "11111111";
  ELSIF (FALLING_EDGE(WR50)) THEN
    DFF_5 <= D;
  END IF;
END PROCESS;

PROCESS(WR51, RESET_n)
BEGIN
  IF (RESET_n = '0') THEN
    DFF_D <= "1111";
    SET_5 <= "1111";
  ELSIF (FALLING_EDGE(WR51)) THEN
    DFF_D <= D(3 DOWNTO 0);
    SET_5 <= D(7 DOWNTO 4);
  END IF;
END PROCESS;

PROCESS(WR60, RESET_n)
BEGIN
  IF (RESET_n = '0') THEN
    DFF_6 <= "11111111";
  ELSIF (FALLING_EDGE(WR60)) THEN
    DFF_6 <= D;
  END IF;
END PROCESS;

PROCESS(WR61, RESET_n)
BEGIN
  IF (RESET_n = '0') THEN
    DFF_E <= "1111";
    SET_6 <= "1111";
  ELSIF (FALLING_EDGE(WR61)) THEN
    DFF_E <= D(3 DOWNTO 0);
    SET_6 <= D(7 DOWNTO 4);
  END IF;
END PROCESS;

PROCESS(WR70, RESET_n)
BEGIN
  IF (RESET_n = '0') THEN
    DFF_7 <= "11111111";
  ELSIF (FALLING_EDGE(WR70)) THEN
    DFF_7 <= D;
  END IF;
END PROCESS;

PROCESS(WR71, RESET_n)
BEGIN
  IF (RESET_n = '0') THEN
    DFF_F <= "1111";
    SET_7 <= "1111";
  ELSIF (FALLING_EDGE(WR71)) THEN
    DFF_F <= D(3 DOWNTO 0);
    SET_7 <= D(7 DOWNTO 4);
  END IF;
END PROCESS;


WITH A(15 DOWNTO 13) SELECT Q_ALT <=
    DFF_8 & DFF_0 WHEN "000",
    DFF_9 & DFF_1 WHEN "001",
    DFF_A & DFF_2 WHEN "010",
    DFF_B & DFF_3 WHEN "011",
    DFF_C & DFF_4 WHEN "100",
    DFF_D & DFF_5 WHEN "101",
    DFF_E & DFF_6 WHEN "110",
    DFF_F & DFF_7 WHEN "111";


Q   <= Q_ALT;
SET <= SET_7 & SET_6 & SET_5 & SET_4 & SET_3 & SET_2 & SET_1 & SET_0;

END bdf_type;